
MACRO rom_data_insel
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN bit7
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 46.00 31.00 48.00 ;
            RECT 24.00 46.00 26.00 48.00 ;
            RECT 19.00 46.00 21.00 48.00 ;
        END
    END bit7
    PIN bit6
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 40.00 31.00 42.00 ;
            RECT 24.00 40.00 26.00 42.00 ;
            RECT 19.00 40.00 21.00 42.00 ;
        END
    END bit6
    PIN bit0
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 4.00 31.00 6.00 ;
            RECT 24.00 4.00 26.00 6.00 ;
            RECT 19.00 4.00 21.00 6.00 ;
        END
    END bit0
    PIN bit1
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 10.00 31.00 12.00 ;
            RECT 24.00 10.00 26.00 12.00 ;
            RECT 19.00 10.00 21.00 12.00 ;
        END
    END bit1
    PIN bit2
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 16.00 31.00 18.00 ;
            RECT 24.00 16.00 26.00 18.00 ;
            RECT 19.00 16.00 21.00 18.00 ;
        END
    END bit2
    PIN bit3
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 22.00 31.00 24.00 ;
            RECT 24.00 22.00 26.00 24.00 ;
            RECT 19.00 22.00 21.00 24.00 ;
        END
    END bit3
    PIN bit4
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 28.00 31.00 30.00 ;
            RECT 24.00 28.00 26.00 30.00 ;
            RECT 19.00 28.00 21.00 30.00 ;
        END
    END bit4
    PIN bit5
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
        END
    END bit5
    PIN prech
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 -1.00 26.00 1.00 ;
        END
    END prech
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 28.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 49.00 11.00 51.00 ;
        RECT 14.00 -1.00 31.00 51.00 ;
    END
END rom_data_insel


MACRO rom_data_invss
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN bit5
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
        END
    END bit5
    PIN bit4
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 28.00 31.00 30.00 ;
            RECT 24.00 28.00 26.00 30.00 ;
            RECT 19.00 28.00 21.00 30.00 ;
        END
    END bit4
    PIN bit3
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 22.00 31.00 24.00 ;
            RECT 24.00 22.00 26.00 24.00 ;
            RECT 19.00 22.00 21.00 24.00 ;
        END
    END bit3
    PIN bit2
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 16.00 31.00 18.00 ;
            RECT 24.00 16.00 26.00 18.00 ;
            RECT 19.00 16.00 21.00 18.00 ;
        END
    END bit2
    PIN bit1
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 10.00 31.00 12.00 ;
            RECT 24.00 10.00 26.00 12.00 ;
            RECT 19.00 10.00 21.00 12.00 ;
        END
    END bit1
    PIN bit0
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 4.00 31.00 6.00 ;
            RECT 24.00 4.00 26.00 6.00 ;
            RECT 19.00 4.00 21.00 6.00 ;
        END
    END bit0
    PIN bit6
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 40.00 31.00 42.00 ;
            RECT 24.00 40.00 26.00 42.00 ;
            RECT 19.00 40.00 21.00 42.00 ;
        END
    END bit6
    PIN bit7
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 46.00 31.00 48.00 ;
            RECT 24.00 46.00 26.00 48.00 ;
            RECT 19.00 46.00 21.00 48.00 ;
        END
    END bit7
    PIN prech
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 49.00 26.00 51.00 ;
        END
    END prech
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 28.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 49.00 11.00 51.00 ;
        RECT 14.00 -1.00 31.00 51.00 ;
    END
END rom_data_invss


MACRO rom_data_midsel
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN bit5
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT -1.00 34.00 1.00 36.00 ;
        END
    END bit5
    PIN bit4
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 28.00 26.00 30.00 ;
            RECT 19.00 28.00 21.00 30.00 ;
            RECT 14.00 28.00 16.00 30.00 ;
            RECT 9.00 28.00 11.00 30.00 ;
            RECT 4.00 28.00 6.00 30.00 ;
            RECT -1.00 28.00 1.00 30.00 ;
        END
    END bit4
    PIN bit3
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 22.00 26.00 24.00 ;
            RECT 19.00 22.00 21.00 24.00 ;
            RECT 14.00 22.00 16.00 24.00 ;
            RECT 9.00 22.00 11.00 24.00 ;
            RECT 4.00 22.00 6.00 24.00 ;
            RECT -1.00 22.00 1.00 24.00 ;
        END
    END bit3
    PIN bit0
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 4.00 26.00 6.00 ;
            RECT 19.00 4.00 21.00 6.00 ;
            RECT 14.00 4.00 16.00 6.00 ;
            RECT 9.00 4.00 11.00 6.00 ;
            RECT 4.00 4.00 6.00 6.00 ;
            RECT -1.00 4.00 1.00 6.00 ;
        END
    END bit0
    PIN bit1
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 10.00 26.00 12.00 ;
            RECT 19.00 10.00 21.00 12.00 ;
            RECT 14.00 10.00 16.00 12.00 ;
            RECT 9.00 10.00 11.00 12.00 ;
            RECT 4.00 10.00 6.00 12.00 ;
            RECT -1.00 10.00 1.00 12.00 ;
        END
    END bit1
    PIN bit2
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 16.00 26.00 18.00 ;
            RECT 19.00 16.00 21.00 18.00 ;
            RECT 14.00 16.00 16.00 18.00 ;
            RECT 9.00 16.00 11.00 18.00 ;
            RECT 4.00 16.00 6.00 18.00 ;
            RECT -1.00 16.00 1.00 18.00 ;
        END
    END bit2
    PIN bit6
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 40.00 26.00 42.00 ;
            RECT 19.00 40.00 21.00 42.00 ;
            RECT 14.00 40.00 16.00 42.00 ;
            RECT 9.00 40.00 11.00 42.00 ;
            RECT 4.00 40.00 6.00 42.00 ;
            RECT -1.00 40.00 1.00 42.00 ;
        END
    END bit6
    PIN bit7
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 46.00 26.00 48.00 ;
            RECT 19.00 46.00 21.00 48.00 ;
            RECT 14.00 46.00 16.00 48.00 ;
            RECT 9.00 46.00 11.00 48.00 ;
            RECT 4.00 46.00 6.00 48.00 ;
            RECT -1.00 46.00 1.00 48.00 ;
        END
    END bit7
    PIN seld
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 -1.00 21.00 1.00 ;
        END
    END seld
    PIN selc
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 -1.00 16.00 1.00 ;
        END
    END selc
    PIN selb
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 -1.00 11.00 1.00 ;
        END
    END selb
    PIN sela
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 -1.00 6.00 1.00 ;
        END
    END sela
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 23.50 48.50 ;
        LAYER L_ALU2 ;
        RECT -1.00 -1.00 26.00 51.00 ;
    END
END rom_data_midsel


MACRO rom_data_midvss
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN bit5
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT -1.00 34.00 1.00 36.00 ;
        END
    END bit5
    PIN bit4
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 28.00 26.00 30.00 ;
            RECT 19.00 28.00 21.00 30.00 ;
            RECT 14.00 28.00 16.00 30.00 ;
            RECT 9.00 28.00 11.00 30.00 ;
            RECT 4.00 28.00 6.00 30.00 ;
            RECT -1.00 28.00 1.00 30.00 ;
        END
    END bit4
    PIN bit3
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 22.00 26.00 24.00 ;
            RECT 19.00 22.00 21.00 24.00 ;
            RECT 14.00 22.00 16.00 24.00 ;
            RECT 9.00 22.00 11.00 24.00 ;
            RECT 4.00 22.00 6.00 24.00 ;
            RECT -1.00 22.00 1.00 24.00 ;
        END
    END bit3
    PIN bit0
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 4.00 26.00 6.00 ;
            RECT 19.00 4.00 21.00 6.00 ;
            RECT 14.00 4.00 16.00 6.00 ;
            RECT 9.00 4.00 11.00 6.00 ;
            RECT 4.00 4.00 6.00 6.00 ;
            RECT -1.00 4.00 1.00 6.00 ;
        END
    END bit0
    PIN bit1
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 10.00 26.00 12.00 ;
            RECT 19.00 10.00 21.00 12.00 ;
            RECT 14.00 10.00 16.00 12.00 ;
            RECT 9.00 10.00 11.00 12.00 ;
            RECT 4.00 10.00 6.00 12.00 ;
            RECT -1.00 10.00 1.00 12.00 ;
        END
    END bit1
    PIN bit2
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 16.00 26.00 18.00 ;
            RECT 19.00 16.00 21.00 18.00 ;
            RECT 14.00 16.00 16.00 18.00 ;
            RECT 9.00 16.00 11.00 18.00 ;
            RECT 4.00 16.00 6.00 18.00 ;
            RECT -1.00 16.00 1.00 18.00 ;
        END
    END bit2
    PIN bit6
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 40.00 26.00 42.00 ;
            RECT 19.00 40.00 21.00 42.00 ;
            RECT 14.00 40.00 16.00 42.00 ;
            RECT 9.00 40.00 11.00 42.00 ;
            RECT 4.00 40.00 6.00 42.00 ;
            RECT -1.00 40.00 1.00 42.00 ;
        END
    END bit6
    PIN bit7
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 46.00 26.00 48.00 ;
            RECT 19.00 46.00 21.00 48.00 ;
            RECT 14.00 46.00 16.00 48.00 ;
            RECT 9.00 46.00 11.00 48.00 ;
            RECT 4.00 46.00 6.00 48.00 ;
            RECT -1.00 46.00 1.00 48.00 ;
        END
    END bit7
    PIN seld
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 49.00 21.00 51.00 ;
        END
    END seld
    PIN selc
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 49.00 16.00 51.00 ;
        END
    END selc
    PIN selb
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 49.00 11.00 51.00 ;
        END
    END selb
    PIN sela
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 49.00 6.00 51.00 ;
        END
    END sela
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 23.50 48.50 ;
        LAYER L_ALU2 ;
        RECT -1.00 -1.00 26.00 51.00 ;
    END
END rom_data_midvss


MACRO rom_data_outsel
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      120.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            LAYER L_ALU3 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
            RECT 109.00 24.00 111.00 26.00 ;
            RECT 109.00 19.00 111.00 21.00 ;
            RECT 109.00 14.00 111.00 16.00 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 109.00 4.00 111.00 6.00 ;
        END
    END q
    PIN bit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 59.00 10.00 61.00 12.00 ;
            RECT 54.00 10.00 56.00 12.00 ;
            RECT 49.00 10.00 51.00 12.00 ;
            RECT 44.00 10.00 46.00 12.00 ;
            RECT 39.00 10.00 41.00 12.00 ;
            RECT 34.00 10.00 36.00 12.00 ;
            RECT 29.00 10.00 31.00 12.00 ;
            RECT 24.00 10.00 26.00 12.00 ;
            RECT 19.00 10.00 21.00 12.00 ;
            RECT 14.00 10.00 16.00 12.00 ;
            RECT 9.00 10.00 11.00 12.00 ;
            RECT 4.00 10.00 6.00 12.00 ;
            RECT -1.00 10.00 1.00 12.00 ;
        END
    END bit1
    PIN bit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 79.00 4.00 81.00 6.00 ;
            RECT 74.00 4.00 76.00 6.00 ;
            RECT 69.00 4.00 71.00 6.00 ;
            RECT 64.00 4.00 66.00 6.00 ;
            RECT 59.00 4.00 61.00 6.00 ;
            RECT 54.00 4.00 56.00 6.00 ;
            RECT 49.00 4.00 51.00 6.00 ;
            RECT 44.00 4.00 46.00 6.00 ;
            RECT 39.00 4.00 41.00 6.00 ;
            RECT 34.00 4.00 36.00 6.00 ;
            RECT 29.00 4.00 31.00 6.00 ;
            RECT 24.00 4.00 26.00 6.00 ;
            RECT 19.00 4.00 21.00 6.00 ;
            RECT 14.00 4.00 16.00 6.00 ;
            RECT 9.00 4.00 11.00 6.00 ;
            RECT 4.00 4.00 6.00 6.00 ;
            RECT -1.00 4.00 1.00 6.00 ;
        END
    END bit0
    PIN bit2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 16.00 41.00 18.00 ;
            RECT 34.00 16.00 36.00 18.00 ;
            RECT 29.00 16.00 31.00 18.00 ;
            RECT 24.00 16.00 26.00 18.00 ;
            RECT 19.00 16.00 21.00 18.00 ;
            RECT 14.00 16.00 16.00 18.00 ;
            RECT 9.00 16.00 11.00 18.00 ;
            RECT 4.00 16.00 6.00 18.00 ;
            RECT -1.00 16.00 1.00 18.00 ;
        END
    END bit2
    PIN bit3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 22.00 21.00 24.00 ;
            RECT 14.00 22.00 16.00 24.00 ;
            RECT 9.00 22.00 11.00 24.00 ;
            RECT 4.00 22.00 6.00 24.00 ;
            RECT -1.00 22.00 1.00 24.00 ;
        END
    END bit3
    PIN bit4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 69.00 28.00 71.00 30.00 ;
            RECT 64.00 28.00 66.00 30.00 ;
            RECT 59.00 28.00 61.00 30.00 ;
            RECT 54.00 28.00 56.00 30.00 ;
            RECT 49.00 28.00 51.00 30.00 ;
            RECT 44.00 28.00 46.00 30.00 ;
            RECT 39.00 28.00 41.00 30.00 ;
            RECT 34.00 28.00 36.00 30.00 ;
            RECT 29.00 28.00 31.00 30.00 ;
            RECT 24.00 28.00 26.00 30.00 ;
            RECT 19.00 28.00 21.00 30.00 ;
            RECT 14.00 28.00 16.00 30.00 ;
            RECT 9.00 28.00 11.00 30.00 ;
            RECT 4.00 28.00 6.00 30.00 ;
            RECT -1.00 28.00 1.00 30.00 ;
        END
    END bit4
    PIN bit7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 46.00 11.00 48.00 ;
            RECT 4.00 46.00 6.00 48.00 ;
            RECT -1.00 46.00 1.00 48.00 ;
        END
    END bit7
    PIN bit5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT -1.00 34.00 1.00 36.00 ;
        END
    END bit5
    PIN bit6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 40.00 31.00 42.00 ;
            RECT 24.00 40.00 26.00 42.00 ;
            RECT 19.00 40.00 21.00 42.00 ;
            RECT 14.00 40.00 16.00 42.00 ;
            RECT 9.00 40.00 11.00 42.00 ;
            RECT 4.00 40.00 6.00 42.00 ;
            RECT -1.00 40.00 1.00 42.00 ;
        END
    END bit6
    PIN mux7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 -1.00 16.00 1.00 ;
        END
    END mux7
    PIN mux3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 -1.00 26.00 1.00 ;
        END
    END mux3
    PIN mux6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 -1.00 36.00 1.00 ;
        END
    END mux6
    PIN mux2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 -1.00 46.00 1.00 ;
        END
    END mux2
    PIN mux5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 54.00 -1.00 56.00 1.00 ;
        END
    END mux5
    PIN mux1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 -1.00 66.00 1.00 ;
        END
    END mux1
    PIN mux4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 74.00 -1.00 76.00 1.00 ;
        END
    END mux4
    PIN mux0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 -1.00 86.00 1.00 ;
        END
    END mux0
    PIN nprech
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 24.00 101.00 26.00 ;
        END
    END nprech
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 118.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 84.00 -1.00 96.00 1.00 ;
        RECT -1.00 -1.00 86.00 51.00 ;
        RECT 84.00 24.00 101.00 26.00 ;
        RECT 84.00 19.00 121.00 21.00 ;
        RECT 84.00 39.00 121.00 41.00 ;
        RECT 93.00 39.00 118.00 41.00 ;
        RECT 87.00 19.00 113.00 21.00 ;
    END
END rom_data_outsel


MACRO rom_data_outsel_ts
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      140.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 124.00 34.00 126.00 36.00 ;
            RECT 119.00 34.00 121.00 36.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            LAYER L_ALU2 ;
            RECT 129.00 9.00 131.00 11.00 ;
            RECT 124.00 9.00 126.00 11.00 ;
            RECT 119.00 9.00 121.00 11.00 ;
            RECT 114.00 9.00 116.00 11.00 ;
            LAYER L_ALU3 ;
            RECT 129.00 44.00 131.00 46.00 ;
            RECT 129.00 39.00 131.00 41.00 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 129.00 29.00 131.00 31.00 ;
            RECT 129.00 24.00 131.00 26.00 ;
            RECT 129.00 19.00 131.00 21.00 ;
            RECT 129.00 14.00 131.00 16.00 ;
            RECT 129.00 9.00 131.00 11.00 ;
            RECT 129.00 4.00 131.00 6.00 ;
        END
    END q
    PIN enx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 24.00 111.00 26.00 ;
        END
    END enx
    PIN nenx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 119.00 24.00 121.00 26.00 ;
        END
    END nenx
    PIN bit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 79.00 4.00 81.00 6.00 ;
            RECT 74.00 4.00 76.00 6.00 ;
            RECT 69.00 4.00 71.00 6.00 ;
            RECT 64.00 4.00 66.00 6.00 ;
            RECT 59.00 4.00 61.00 6.00 ;
            RECT 54.00 4.00 56.00 6.00 ;
            RECT 49.00 4.00 51.00 6.00 ;
            RECT 44.00 4.00 46.00 6.00 ;
            RECT 39.00 4.00 41.00 6.00 ;
            RECT 34.00 4.00 36.00 6.00 ;
            RECT 29.00 4.00 31.00 6.00 ;
            RECT 24.00 4.00 26.00 6.00 ;
            RECT 19.00 4.00 21.00 6.00 ;
            RECT 14.00 4.00 16.00 6.00 ;
            RECT 9.00 4.00 11.00 6.00 ;
            RECT 4.00 4.00 6.00 6.00 ;
            RECT -1.00 4.00 1.00 6.00 ;
        END
    END bit0
    PIN bit2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 16.00 41.00 18.00 ;
            RECT 34.00 16.00 36.00 18.00 ;
            RECT 29.00 16.00 31.00 18.00 ;
            RECT 24.00 16.00 26.00 18.00 ;
            RECT 19.00 16.00 21.00 18.00 ;
            RECT 14.00 16.00 16.00 18.00 ;
            RECT 9.00 16.00 11.00 18.00 ;
            RECT 4.00 16.00 6.00 18.00 ;
            RECT -1.00 16.00 1.00 18.00 ;
        END
    END bit2
    PIN bit3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 22.00 21.00 24.00 ;
            RECT 14.00 22.00 16.00 24.00 ;
            RECT 9.00 22.00 11.00 24.00 ;
            RECT 4.00 22.00 6.00 24.00 ;
            RECT -1.00 22.00 1.00 24.00 ;
        END
    END bit3
    PIN bit4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 69.00 28.00 71.00 30.00 ;
            RECT 64.00 28.00 66.00 30.00 ;
            RECT 59.00 28.00 61.00 30.00 ;
            RECT 54.00 28.00 56.00 30.00 ;
            RECT 49.00 28.00 51.00 30.00 ;
            RECT 44.00 28.00 46.00 30.00 ;
            RECT 39.00 28.00 41.00 30.00 ;
            RECT 34.00 28.00 36.00 30.00 ;
            RECT 29.00 28.00 31.00 30.00 ;
            RECT 24.00 28.00 26.00 30.00 ;
            RECT 19.00 28.00 21.00 30.00 ;
            RECT 14.00 28.00 16.00 30.00 ;
            RECT 9.00 28.00 11.00 30.00 ;
            RECT 4.00 28.00 6.00 30.00 ;
            RECT -1.00 28.00 1.00 30.00 ;
        END
    END bit4
    PIN bit7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 46.00 11.00 48.00 ;
            RECT 4.00 46.00 6.00 48.00 ;
            RECT -1.00 46.00 1.00 48.00 ;
        END
    END bit7
    PIN bit5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT -1.00 34.00 1.00 36.00 ;
        END
    END bit5
    PIN bit6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 40.00 31.00 42.00 ;
            RECT 24.00 40.00 26.00 42.00 ;
            RECT 19.00 40.00 21.00 42.00 ;
            RECT 14.00 40.00 16.00 42.00 ;
            RECT 9.00 40.00 11.00 42.00 ;
            RECT 4.00 40.00 6.00 42.00 ;
            RECT -1.00 40.00 1.00 42.00 ;
        END
    END bit6
    PIN mux7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 -1.00 16.00 1.00 ;
        END
    END mux7
    PIN mux3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 -1.00 26.00 1.00 ;
        END
    END mux3
    PIN mux6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 -1.00 36.00 1.00 ;
        END
    END mux6
    PIN mux2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 -1.00 46.00 1.00 ;
        END
    END mux2
    PIN mux5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 54.00 -1.00 56.00 1.00 ;
        END
    END mux5
    PIN mux1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 -1.00 66.00 1.00 ;
        END
    END mux1
    PIN mux4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 74.00 -1.00 76.00 1.00 ;
        END
    END mux4
    PIN mux0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 -1.00 86.00 1.00 ;
        END
    END mux0
    PIN nprech
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 24.00 101.00 26.00 ;
        END
    END nprech
    PIN bit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 59.00 10.00 61.00 12.00 ;
            RECT 54.00 10.00 56.00 12.00 ;
            RECT 49.00 10.00 51.00 12.00 ;
            RECT 44.00 10.00 46.00 12.00 ;
            RECT 39.00 10.00 41.00 12.00 ;
            RECT 34.00 10.00 36.00 12.00 ;
            RECT 29.00 10.00 31.00 12.00 ;
            RECT 24.00 10.00 26.00 12.00 ;
            RECT 19.00 10.00 21.00 12.00 ;
            RECT 14.00 10.00 16.00 12.00 ;
            RECT 9.00 10.00 11.00 12.00 ;
            RECT 4.00 10.00 6.00 12.00 ;
            RECT -1.00 10.00 1.00 12.00 ;
        END
    END bit1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 138.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 84.00 14.00 121.00 16.00 ;
        RECT 87.00 14.00 121.00 16.00 ;
        RECT 93.00 39.00 134.00 41.00 ;
        RECT -1.00 -1.00 86.00 51.00 ;
        RECT 84.00 39.00 136.00 41.00 ;
        RECT 84.00 24.00 121.00 26.00 ;
    END
END rom_data_outsel_ts


MACRO rom_data_outvss
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      120.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
            RECT 109.00 24.00 111.00 26.00 ;
            RECT 109.00 19.00 111.00 21.00 ;
            RECT 109.00 14.00 111.00 16.00 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 109.00 4.00 111.00 6.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
        END
    END q
    PIN nprech
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 24.00 101.00 26.00 ;
        END
    END nprech
    PIN bit6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 40.00 31.00 42.00 ;
            RECT 24.00 40.00 26.00 42.00 ;
            RECT 19.00 40.00 21.00 42.00 ;
            RECT 14.00 40.00 16.00 42.00 ;
            RECT 9.00 40.00 11.00 42.00 ;
            RECT 4.00 40.00 6.00 42.00 ;
            RECT -1.00 40.00 1.00 42.00 ;
        END
    END bit6
    PIN bit5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT -1.00 34.00 1.00 36.00 ;
        END
    END bit5
    PIN bit7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 46.00 11.00 48.00 ;
            RECT 4.00 46.00 6.00 48.00 ;
            RECT -1.00 46.00 1.00 48.00 ;
        END
    END bit7
    PIN bit4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 69.00 28.00 71.00 30.00 ;
            RECT 64.00 28.00 66.00 30.00 ;
            RECT 59.00 28.00 61.00 30.00 ;
            RECT 54.00 28.00 56.00 30.00 ;
            RECT 49.00 28.00 51.00 30.00 ;
            RECT 44.00 28.00 46.00 30.00 ;
            RECT 39.00 28.00 41.00 30.00 ;
            RECT 34.00 28.00 36.00 30.00 ;
            RECT 29.00 28.00 31.00 30.00 ;
            RECT 24.00 28.00 26.00 30.00 ;
            RECT 19.00 28.00 21.00 30.00 ;
            RECT 14.00 28.00 16.00 30.00 ;
            RECT 9.00 28.00 11.00 30.00 ;
            RECT 4.00 28.00 6.00 30.00 ;
            RECT -1.00 28.00 1.00 30.00 ;
        END
    END bit4
    PIN bit3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 22.00 21.00 24.00 ;
            RECT 14.00 22.00 16.00 24.00 ;
            RECT 9.00 22.00 11.00 24.00 ;
            RECT 4.00 22.00 6.00 24.00 ;
            RECT -1.00 22.00 1.00 24.00 ;
        END
    END bit3
    PIN bit2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 16.00 41.00 18.00 ;
            RECT 34.00 16.00 36.00 18.00 ;
            RECT 29.00 16.00 31.00 18.00 ;
            RECT 24.00 16.00 26.00 18.00 ;
            RECT 19.00 16.00 21.00 18.00 ;
            RECT 14.00 16.00 16.00 18.00 ;
            RECT 9.00 16.00 11.00 18.00 ;
            RECT 4.00 16.00 6.00 18.00 ;
            RECT -1.00 16.00 1.00 18.00 ;
        END
    END bit2
    PIN bit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 79.00 4.00 81.00 6.00 ;
            RECT 74.00 4.00 76.00 6.00 ;
            RECT 69.00 4.00 71.00 6.00 ;
            RECT 64.00 4.00 66.00 6.00 ;
            RECT 59.00 4.00 61.00 6.00 ;
            RECT 54.00 4.00 56.00 6.00 ;
            RECT 49.00 4.00 51.00 6.00 ;
            RECT 44.00 4.00 46.00 6.00 ;
            RECT 39.00 4.00 41.00 6.00 ;
            RECT 34.00 4.00 36.00 6.00 ;
            RECT 29.00 4.00 31.00 6.00 ;
            RECT 24.00 4.00 26.00 6.00 ;
            RECT 19.00 4.00 21.00 6.00 ;
            RECT 14.00 4.00 16.00 6.00 ;
            RECT 9.00 4.00 11.00 6.00 ;
            RECT 4.00 4.00 6.00 6.00 ;
            RECT -1.00 4.00 1.00 6.00 ;
        END
    END bit0
    PIN mux0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 49.00 86.00 51.00 ;
        END
    END mux0
    PIN mux4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 74.00 49.00 76.00 51.00 ;
        END
    END mux4
    PIN mux1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 49.00 66.00 51.00 ;
        END
    END mux1
    PIN mux5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 54.00 49.00 56.00 51.00 ;
        END
    END mux5
    PIN mux2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 49.00 46.00 51.00 ;
        END
    END mux2
    PIN mux6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 49.00 36.00 51.00 ;
        END
    END mux6
    PIN mux3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 49.00 26.00 51.00 ;
        END
    END mux3
    PIN mux7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 49.00 16.00 51.00 ;
        END
    END mux7
    PIN bit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 59.00 10.00 61.00 12.00 ;
            RECT 54.00 10.00 56.00 12.00 ;
            RECT 49.00 10.00 51.00 12.00 ;
            RECT 44.00 10.00 46.00 12.00 ;
            RECT 39.00 10.00 41.00 12.00 ;
            RECT 34.00 10.00 36.00 12.00 ;
            RECT 29.00 10.00 31.00 12.00 ;
            RECT 24.00 10.00 26.00 12.00 ;
            RECT 19.00 10.00 21.00 12.00 ;
            RECT 14.00 10.00 16.00 12.00 ;
            RECT 9.00 10.00 11.00 12.00 ;
            RECT 4.00 10.00 6.00 12.00 ;
            RECT -1.00 10.00 1.00 12.00 ;
        END
    END bit1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 118.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 84.00 24.00 101.00 26.00 ;
        RECT 87.00 19.00 113.00 21.00 ;
        RECT 93.00 39.00 118.00 41.00 ;
        RECT -1.00 -1.00 86.00 51.00 ;
        RECT 84.00 39.00 121.00 41.00 ;
        RECT 84.00 19.00 121.00 21.00 ;
    END
END rom_data_outvss


MACRO rom_data_outvss_ts
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      140.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU3 ;
            RECT 129.00 44.00 131.00 46.00 ;
            RECT 129.00 39.00 131.00 41.00 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 129.00 29.00 131.00 31.00 ;
            RECT 129.00 24.00 131.00 26.00 ;
            RECT 129.00 19.00 131.00 21.00 ;
            RECT 129.00 14.00 131.00 16.00 ;
            RECT 129.00 9.00 131.00 11.00 ;
            RECT 129.00 4.00 131.00 6.00 ;
            LAYER L_ALU2 ;
            RECT 129.00 9.00 131.00 11.00 ;
            RECT 124.00 9.00 126.00 11.00 ;
            RECT 119.00 9.00 121.00 11.00 ;
            RECT 114.00 9.00 116.00 11.00 ;
            LAYER L_ALU2 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 124.00 34.00 126.00 36.00 ;
            RECT 119.00 34.00 121.00 36.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
        END
    END q
    PIN mux0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 49.00 86.00 51.00 ;
        END
    END mux0
    PIN mux4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 74.00 49.00 76.00 51.00 ;
        END
    END mux4
    PIN mux1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 49.00 66.00 51.00 ;
        END
    END mux1
    PIN mux5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 54.00 49.00 56.00 51.00 ;
        END
    END mux5
    PIN mux2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 49.00 46.00 51.00 ;
        END
    END mux2
    PIN mux6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 49.00 36.00 51.00 ;
        END
    END mux6
    PIN mux3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 49.00 26.00 51.00 ;
        END
    END mux3
    PIN mux7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 49.00 16.00 51.00 ;
        END
    END mux7
    PIN nprech
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 24.00 101.00 26.00 ;
        END
    END nprech
    PIN bit6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 40.00 31.00 42.00 ;
            RECT 24.00 40.00 26.00 42.00 ;
            RECT 19.00 40.00 21.00 42.00 ;
            RECT 14.00 40.00 16.00 42.00 ;
            RECT 9.00 40.00 11.00 42.00 ;
            RECT 4.00 40.00 6.00 42.00 ;
            RECT -1.00 40.00 1.00 42.00 ;
        END
    END bit6
    PIN bit5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT -1.00 34.00 1.00 36.00 ;
        END
    END bit5
    PIN bit7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 46.00 11.00 48.00 ;
            RECT 4.00 46.00 6.00 48.00 ;
            RECT -1.00 46.00 1.00 48.00 ;
        END
    END bit7
    PIN bit4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 69.00 28.00 71.00 30.00 ;
            RECT 64.00 28.00 66.00 30.00 ;
            RECT 59.00 28.00 61.00 30.00 ;
            RECT 54.00 28.00 56.00 30.00 ;
            RECT 49.00 28.00 51.00 30.00 ;
            RECT 44.00 28.00 46.00 30.00 ;
            RECT 39.00 28.00 41.00 30.00 ;
            RECT 34.00 28.00 36.00 30.00 ;
            RECT 29.00 28.00 31.00 30.00 ;
            RECT 24.00 28.00 26.00 30.00 ;
            RECT 19.00 28.00 21.00 30.00 ;
            RECT 14.00 28.00 16.00 30.00 ;
            RECT 9.00 28.00 11.00 30.00 ;
            RECT 4.00 28.00 6.00 30.00 ;
            RECT -1.00 28.00 1.00 30.00 ;
        END
    END bit4
    PIN bit3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 22.00 21.00 24.00 ;
            RECT 14.00 22.00 16.00 24.00 ;
            RECT 9.00 22.00 11.00 24.00 ;
            RECT 4.00 22.00 6.00 24.00 ;
            RECT -1.00 22.00 1.00 24.00 ;
        END
    END bit3
    PIN bit2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 16.00 41.00 18.00 ;
            RECT 34.00 16.00 36.00 18.00 ;
            RECT 29.00 16.00 31.00 18.00 ;
            RECT 24.00 16.00 26.00 18.00 ;
            RECT 19.00 16.00 21.00 18.00 ;
            RECT 14.00 16.00 16.00 18.00 ;
            RECT 9.00 16.00 11.00 18.00 ;
            RECT 4.00 16.00 6.00 18.00 ;
            RECT -1.00 16.00 1.00 18.00 ;
        END
    END bit2
    PIN bit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 79.00 4.00 81.00 6.00 ;
            RECT 74.00 4.00 76.00 6.00 ;
            RECT 69.00 4.00 71.00 6.00 ;
            RECT 64.00 4.00 66.00 6.00 ;
            RECT 59.00 4.00 61.00 6.00 ;
            RECT 54.00 4.00 56.00 6.00 ;
            RECT 49.00 4.00 51.00 6.00 ;
            RECT 44.00 4.00 46.00 6.00 ;
            RECT 39.00 4.00 41.00 6.00 ;
            RECT 34.00 4.00 36.00 6.00 ;
            RECT 29.00 4.00 31.00 6.00 ;
            RECT 24.00 4.00 26.00 6.00 ;
            RECT 19.00 4.00 21.00 6.00 ;
            RECT 14.00 4.00 16.00 6.00 ;
            RECT 9.00 4.00 11.00 6.00 ;
            RECT 4.00 4.00 6.00 6.00 ;
            RECT -1.00 4.00 1.00 6.00 ;
        END
    END bit0
    PIN nenx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 119.00 24.00 121.00 26.00 ;
        END
    END nenx
    PIN enx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 24.00 111.00 26.00 ;
        END
    END enx
    PIN bit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 59.00 10.00 61.00 12.00 ;
            RECT 54.00 10.00 56.00 12.00 ;
            RECT 49.00 10.00 51.00 12.00 ;
            RECT 44.00 10.00 46.00 12.00 ;
            RECT 39.00 10.00 41.00 12.00 ;
            RECT 34.00 10.00 36.00 12.00 ;
            RECT 29.00 10.00 31.00 12.00 ;
            RECT 24.00 10.00 26.00 12.00 ;
            RECT 19.00 10.00 21.00 12.00 ;
            RECT 14.00 10.00 16.00 12.00 ;
            RECT 9.00 10.00 11.00 12.00 ;
            RECT 4.00 10.00 6.00 12.00 ;
            RECT -1.00 10.00 1.00 12.00 ;
        END
    END bit1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 138.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 84.00 24.00 121.00 26.00 ;
        RECT 84.00 39.00 136.00 41.00 ;
        RECT 84.00 14.00 121.00 16.00 ;
        RECT 93.00 39.00 134.00 41.00 ;
        RECT -1.00 -1.00 86.00 51.00 ;
        RECT 87.00 14.00 121.00 16.00 ;
    END
END rom_data_outvss_ts


MACRO rom_dec_adbuf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nadx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 34.00 11.00 36.00 ;
        END
    END nadx
    PIN adx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 44.00 26.00 46.00 ;
        END
    END adx
    PIN ad
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END ad
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 28.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 9.00 39.00 26.00 41.00 ;
        RECT 20.00 39.00 26.00 41.00 ;
        RECT 24.00 39.00 26.00 46.00 ;
    END
END rom_dec_adbuf


MACRO rom_dec_col2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 29.00 31.00 31.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 29.00 11.00 31.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END i0
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 48.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 29.00 31.00 31.00 ;
    END
END rom_dec_col2


MACRO rom_dec_col3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 29.00 31.00 31.00 ;
        END
    END q
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 29.00 21.00 31.00 ;
        END
    END i2
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 29.00 11.00 31.00 ;
        END
    END i1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 48.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 29.00 31.00 31.00 ;
    END
END rom_dec_col3


MACRO rom_dec_col4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 29.00 31.00 31.00 ;
        END
    END q
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 29.00 21.00 31.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 29.00 16.00 31.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 29.00 11.00 31.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END i0
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 48.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 29.00 29.00 41.00 31.00 ;
        RECT 4.00 29.00 41.00 31.00 ;
        RECT 19.00 29.00 23.00 31.00 ;
    END
END rom_dec_col4


MACRO rom_dec_colbuf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nax
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 29.00 21.00 31.00 ;
        END
    END nax
    PIN ax
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 29.00 11.00 31.00 ;
        END
    END ax
    PIN a
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 29.00 16.00 31.00 ;
        END
    END a
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 28.50 48.50 ;
        LAYER L_ALU2 ;
        RECT 9.00 29.00 21.00 31.00 ;
    END
END rom_dec_colbuf


MACRO rom_dec_line01
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN col
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
        END
    END col
    PIN nck0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nck0
    PIN nck1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 89.00 41.00 91.00 ;
        END
    END nck1
    PIN sel1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 84.00 36.00 86.00 ;
        END
    END sel1
    PIN sel0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END sel0
    PIN line1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END line1
    PIN line0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 79.00 6.00 81.00 ;
        END
    END line0
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 48.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 24.00 31.00 26.00 ;
        RECT -1.00 19.00 51.00 21.00 ;
        RECT -1.00 24.00 51.00 26.00 ;
        RECT -1.00 79.00 51.00 81.00 ;
        RECT -1.00 74.00 51.00 76.00 ;
    END
END rom_dec_line01


MACRO rom_dec_line23
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN col
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
        END
    END col
    PIN line3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END line3
    PIN line2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 79.00 11.00 81.00 ;
        END
    END line2
    PIN nck2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nck2
    PIN sel2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END sel2
    PIN sel3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 84.00 36.00 86.00 ;
        END
    END sel3
    PIN nck3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 89.00 41.00 91.00 ;
        END
    END nck3
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 48.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 24.00 31.00 26.00 ;
        RECT -1.00 79.00 51.00 81.00 ;
        RECT -1.00 74.00 51.00 76.00 ;
        RECT -1.00 19.00 51.00 21.00 ;
        RECT -1.00 24.00 51.00 26.00 ;
    END
END rom_dec_line23


MACRO rom_dec_line45
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN col
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
        END
    END col
    PIN nck4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nck4
    PIN nck5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 89.00 41.00 91.00 ;
        END
    END nck5
    PIN sel4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END sel4
    PIN sel5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 84.00 36.00 86.00 ;
        END
    END sel5
    PIN line4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 79.00 16.00 81.00 ;
        END
    END line4
    PIN line5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END line5
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 48.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 24.00 31.00 26.00 ;
        RECT -1.00 19.00 51.00 21.00 ;
        RECT -1.00 24.00 51.00 26.00 ;
        RECT -1.00 74.00 51.00 76.00 ;
        RECT -1.00 79.00 51.00 81.00 ;
    END
END rom_dec_line45


MACRO rom_dec_line67
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN col
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
        END
    END col
    PIN nck6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nck6
    PIN nck7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 89.00 41.00 91.00 ;
        END
    END nck7
    PIN sel6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END sel6
    PIN sel7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 84.00 36.00 86.00 ;
        END
    END sel7
    PIN line6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 79.00 21.00 81.00 ;
        END
    END line6
    PIN line7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END line7
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 48.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 24.00 31.00 26.00 ;
        RECT -1.00 19.00 51.00 21.00 ;
        RECT -1.00 24.00 51.00 26.00 ;
        RECT -1.00 74.00 51.00 76.00 ;
        RECT -1.00 79.00 51.00 81.00 ;
    END
END rom_dec_line67


MACRO rom_dec_nop
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 28.50 48.50 ;
    END
END rom_dec_nop


MACRO rom_dec_prech
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN nprech
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 14.00 64.00 16.00 66.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
        END
    END nprech
    PIN prech
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 79.00 26.00 81.00 ;
            RECT 24.00 74.00 26.00 76.00 ;
            RECT 24.00 69.00 26.00 71.00 ;
            RECT 24.00 64.00 26.00 66.00 ;
            RECT 24.00 59.00 26.00 61.00 ;
            RECT 24.00 54.00 26.00 56.00 ;
            RECT 24.00 49.00 26.00 51.00 ;
            RECT 24.00 44.00 26.00 46.00 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END prech
    PIN nck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 28.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 14.00 79.00 26.00 81.00 ;
        RECT 4.00 19.00 26.00 21.00 ;
        RECT 8.00 19.00 26.00 21.00 ;
    END
END rom_dec_prech


MACRO rom_dec_selmux01
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      120.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN sel1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel1
    PIN mux1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 59.00 66.00 61.00 ;
        END
    END mux1
    PIN mux0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 39.00 86.00 41.00 ;
        END
    END mux0
    PIN sel0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel0
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 104.00 84.00 106.00 86.00 ;
            RECT 104.00 79.00 106.00 81.00 ;
            RECT 104.00 74.00 106.00 76.00 ;
            RECT 104.00 69.00 106.00 71.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 104.00 59.00 106.00 61.00 ;
            RECT 104.00 54.00 106.00 56.00 ;
            RECT 104.00 49.00 106.00 51.00 ;
            RECT 104.00 44.00 106.00 46.00 ;
            RECT 104.00 39.00 106.00 41.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 104.00 29.00 106.00 31.00 ;
            RECT 104.00 24.00 106.00 26.00 ;
            RECT 104.00 19.00 106.00 21.00 ;
            RECT 104.00 14.00 106.00 16.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
            RECT 84.00 9.00 86.00 11.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
            RECT 74.00 9.00 76.00 11.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
            RECT 64.00 9.00 66.00 11.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 89.00 111.00 91.00 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 84.00 89.00 86.00 91.00 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 4.00 89.00 6.00 91.00 ;
        END
    END nck
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END selrom
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 74.00 116.00 76.00 ;
            RECT 114.00 69.00 116.00 71.00 ;
            RECT 114.00 64.00 116.00 66.00 ;
            RECT 114.00 59.00 116.00 61.00 ;
            RECT 114.00 54.00 116.00 56.00 ;
            RECT 114.00 49.00 116.00 51.00 ;
            RECT 114.00 44.00 116.00 46.00 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
        END
    END ck
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
        END
    END a5
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 118.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 64.00 79.00 96.00 81.00 ;
        RECT 64.00 19.00 96.00 21.00 ;
        RECT 9.00 59.00 66.00 61.00 ;
        RECT 9.00 59.00 66.00 61.00 ;
        RECT 79.00 69.00 111.00 71.00 ;
        RECT 29.00 74.00 41.00 76.00 ;
        RECT 44.00 79.00 51.00 81.00 ;
        RECT 59.00 74.00 91.00 76.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 59.00 24.00 91.00 26.00 ;
        RECT 44.00 19.00 51.00 21.00 ;
        RECT 29.00 24.00 41.00 26.00 ;
        RECT 79.00 29.00 111.00 31.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 9.00 39.00 85.00 41.00 ;
        RECT 4.00 19.00 116.00 21.00 ;
        RECT 4.00 24.00 116.00 26.00 ;
        RECT 4.00 29.00 116.00 31.00 ;
        RECT 4.00 39.00 116.00 41.00 ;
        RECT 4.00 59.00 116.00 61.00 ;
        RECT 4.00 69.00 116.00 71.00 ;
        RECT 4.00 74.00 116.00 76.00 ;
        RECT 4.00 79.00 116.00 81.00 ;
    END
END rom_dec_selmux01


MACRO rom_dec_selmux01_ts
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      140.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN enx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END enx
    PIN nenx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 119.00 74.00 121.00 76.00 ;
            RECT 119.00 69.00 121.00 71.00 ;
            RECT 119.00 64.00 121.00 66.00 ;
            RECT 119.00 59.00 121.00 61.00 ;
            RECT 119.00 54.00 121.00 56.00 ;
            RECT 119.00 49.00 121.00 51.00 ;
            RECT 119.00 44.00 121.00 46.00 ;
            RECT 119.00 39.00 121.00 41.00 ;
            RECT 119.00 34.00 121.00 36.00 ;
            RECT 119.00 29.00 121.00 31.00 ;
            RECT 119.00 24.00 121.00 26.00 ;
        END
    END nenx
    PIN sel1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel1
    PIN mux1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 59.00 66.00 61.00 ;
        END
    END mux1
    PIN mux0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 39.00 86.00 41.00 ;
        END
    END mux0
    PIN sel0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel0
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 104.00 84.00 106.00 86.00 ;
            RECT 104.00 79.00 106.00 81.00 ;
            RECT 104.00 74.00 106.00 76.00 ;
            RECT 104.00 69.00 106.00 71.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 104.00 59.00 106.00 61.00 ;
            RECT 104.00 54.00 106.00 56.00 ;
            RECT 104.00 49.00 106.00 51.00 ;
            RECT 104.00 44.00 106.00 46.00 ;
            RECT 104.00 39.00 106.00 41.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 104.00 29.00 106.00 31.00 ;
            RECT 104.00 24.00 106.00 26.00 ;
            RECT 104.00 19.00 106.00 21.00 ;
            RECT 104.00 14.00 106.00 16.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
            RECT 84.00 9.00 86.00 11.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
            RECT 74.00 9.00 76.00 11.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
            RECT 64.00 9.00 66.00 11.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 89.00 111.00 91.00 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 84.00 89.00 86.00 91.00 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 4.00 89.00 6.00 91.00 ;
        END
    END nck
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 74.00 116.00 76.00 ;
            RECT 114.00 69.00 116.00 71.00 ;
            RECT 114.00 64.00 116.00 66.00 ;
            RECT 114.00 59.00 116.00 61.00 ;
            RECT 114.00 54.00 116.00 56.00 ;
            RECT 114.00 49.00 116.00 51.00 ;
            RECT 114.00 44.00 116.00 46.00 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
        END
    END ck
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 129.00 79.00 131.00 81.00 ;
            RECT 129.00 74.00 131.00 76.00 ;
            RECT 129.00 69.00 131.00 71.00 ;
            RECT 129.00 64.00 131.00 66.00 ;
            RECT 129.00 59.00 131.00 61.00 ;
            RECT 129.00 54.00 131.00 56.00 ;
            RECT 129.00 49.00 131.00 51.00 ;
            RECT 129.00 44.00 131.00 46.00 ;
            RECT 129.00 39.00 131.00 41.00 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 129.00 29.00 131.00 31.00 ;
            RECT 129.00 24.00 131.00 26.00 ;
            RECT 129.00 19.00 131.00 21.00 ;
        END
    END selrom
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
        END
    END a5
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 138.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 119.00 24.00 136.00 26.00 ;
        RECT 119.00 74.00 136.00 76.00 ;
        RECT 4.00 19.00 136.00 21.00 ;
        RECT 4.00 79.00 136.00 81.00 ;
        RECT 64.00 79.00 96.00 81.00 ;
        RECT 64.00 19.00 96.00 21.00 ;
        RECT 9.00 59.00 66.00 61.00 ;
        RECT 29.00 74.00 41.00 76.00 ;
        RECT 44.00 79.00 51.00 81.00 ;
        RECT 59.00 74.00 91.00 76.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 59.00 24.00 91.00 26.00 ;
        RECT 44.00 19.00 51.00 21.00 ;
        RECT 29.00 24.00 41.00 26.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 9.00 39.00 85.00 41.00 ;
        RECT 4.00 24.00 136.00 26.00 ;
        RECT 4.00 39.00 86.00 41.00 ;
        RECT 9.00 59.00 66.00 61.00 ;
        RECT 4.00 74.00 136.00 76.00 ;
        RECT 4.00 59.00 66.00 61.00 ;
        RECT 79.00 29.00 125.00 31.00 ;
        RECT 79.00 69.00 125.00 71.00 ;
        RECT 4.00 69.00 136.00 71.00 ;
        RECT 4.00 29.00 136.00 31.00 ;
    END
END rom_dec_selmux01_ts


MACRO rom_dec_selmux23
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      120.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN sel2
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel2
    PIN sel3
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel3
    PIN mux3
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 59.00 26.00 61.00 ;
        END
    END mux3
    PIN mux2
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 39.00 46.00 41.00 ;
        END
    END mux2
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 104.00 84.00 106.00 86.00 ;
            RECT 104.00 79.00 106.00 81.00 ;
            RECT 104.00 74.00 106.00 76.00 ;
            RECT 104.00 69.00 106.00 71.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 104.00 59.00 106.00 61.00 ;
            RECT 104.00 54.00 106.00 56.00 ;
            RECT 104.00 49.00 106.00 51.00 ;
            RECT 104.00 44.00 106.00 46.00 ;
            RECT 104.00 39.00 106.00 41.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 104.00 29.00 106.00 31.00 ;
            RECT 104.00 24.00 106.00 26.00 ;
            RECT 104.00 19.00 106.00 21.00 ;
            RECT 104.00 14.00 106.00 16.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 89.00 111.00 91.00 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 84.00 89.00 86.00 91.00 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 4.00 89.00 6.00 91.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
            RECT 84.00 9.00 86.00 11.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
            RECT 74.00 9.00 76.00 11.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
            RECT 64.00 9.00 66.00 11.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END nck
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 74.00 116.00 76.00 ;
            RECT 114.00 69.00 116.00 71.00 ;
            RECT 114.00 64.00 116.00 66.00 ;
            RECT 114.00 59.00 116.00 61.00 ;
            RECT 114.00 54.00 116.00 56.00 ;
            RECT 114.00 49.00 116.00 51.00 ;
            RECT 114.00 44.00 116.00 46.00 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
        END
    END ck
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END selrom
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
            RECT 99.00 54.00 101.00 56.00 ;
            RECT 99.00 49.00 101.00 51.00 ;
            RECT 99.00 44.00 101.00 46.00 ;
            RECT 99.00 39.00 101.00 41.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
            RECT 99.00 14.00 101.00 16.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
        END
    END a5
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 118.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 79.00 116.00 81.00 ;
        RECT 4.00 74.00 116.00 76.00 ;
        RECT 4.00 69.00 116.00 71.00 ;
        RECT 4.00 59.00 116.00 61.00 ;
        RECT 4.00 39.00 116.00 41.00 ;
        RECT 4.00 29.00 116.00 31.00 ;
        RECT 4.00 24.00 116.00 26.00 ;
        RECT 4.00 19.00 116.00 21.00 ;
        RECT 64.00 19.00 96.00 21.00 ;
        RECT 64.00 79.00 96.00 81.00 ;
        RECT 19.00 74.00 41.00 76.00 ;
        RECT 59.00 74.00 81.00 76.00 ;
        RECT 59.00 24.00 81.00 26.00 ;
        RECT 19.00 24.00 41.00 26.00 ;
        RECT 9.00 39.00 46.00 41.00 ;
        RECT 9.00 59.00 26.00 61.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 79.00 29.00 111.00 31.00 ;
        RECT 44.00 19.00 51.00 21.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 44.00 79.00 51.00 81.00 ;
        RECT 79.00 69.00 111.00 71.00 ;
    END
END rom_dec_selmux23


MACRO rom_dec_selmux23_ts
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      140.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN mux3
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 59.00 26.00 61.00 ;
        END
    END mux3
    PIN mux2
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 39.00 46.00 41.00 ;
        END
    END mux2
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 109.00 89.00 111.00 91.00 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 84.00 89.00 86.00 91.00 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 4.00 89.00 6.00 91.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
            RECT 84.00 9.00 86.00 11.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
            RECT 74.00 9.00 76.00 11.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
            RECT 64.00 9.00 66.00 11.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
            LAYER L_ALU3 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 104.00 84.00 106.00 86.00 ;
            RECT 104.00 79.00 106.00 81.00 ;
            RECT 104.00 74.00 106.00 76.00 ;
            RECT 104.00 69.00 106.00 71.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 104.00 59.00 106.00 61.00 ;
            RECT 104.00 54.00 106.00 56.00 ;
            RECT 104.00 49.00 106.00 51.00 ;
            RECT 104.00 44.00 106.00 46.00 ;
            RECT 104.00 39.00 106.00 41.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 104.00 29.00 106.00 31.00 ;
            RECT 104.00 24.00 106.00 26.00 ;
            RECT 104.00 19.00 106.00 21.00 ;
            RECT 104.00 14.00 106.00 16.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
        END
    END nck
    PIN sel2
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel2
    PIN sel3
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel3
    PIN enx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END enx
    PIN nenx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 119.00 74.00 121.00 76.00 ;
            RECT 119.00 69.00 121.00 71.00 ;
            RECT 119.00 64.00 121.00 66.00 ;
            RECT 119.00 59.00 121.00 61.00 ;
            RECT 119.00 54.00 121.00 56.00 ;
            RECT 119.00 49.00 121.00 51.00 ;
            RECT 119.00 44.00 121.00 46.00 ;
            RECT 119.00 39.00 121.00 41.00 ;
            RECT 119.00 34.00 121.00 36.00 ;
            RECT 119.00 29.00 121.00 31.00 ;
            RECT 119.00 24.00 121.00 26.00 ;
        END
    END nenx
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
            RECT 99.00 54.00 101.00 56.00 ;
            RECT 99.00 49.00 101.00 51.00 ;
            RECT 99.00 44.00 101.00 46.00 ;
            RECT 99.00 39.00 101.00 41.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
            RECT 99.00 14.00 101.00 16.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
        END
    END a5
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 74.00 116.00 76.00 ;
            RECT 114.00 69.00 116.00 71.00 ;
            RECT 114.00 64.00 116.00 66.00 ;
            RECT 114.00 59.00 116.00 61.00 ;
            RECT 114.00 54.00 116.00 56.00 ;
            RECT 114.00 49.00 116.00 51.00 ;
            RECT 114.00 44.00 116.00 46.00 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
        END
    END ck
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 129.00 79.00 131.00 81.00 ;
            RECT 129.00 74.00 131.00 76.00 ;
            RECT 129.00 69.00 131.00 71.00 ;
            RECT 129.00 64.00 131.00 66.00 ;
            RECT 129.00 59.00 131.00 61.00 ;
            RECT 129.00 54.00 131.00 56.00 ;
            RECT 129.00 49.00 131.00 51.00 ;
            RECT 129.00 44.00 131.00 46.00 ;
            RECT 129.00 39.00 131.00 41.00 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 129.00 29.00 131.00 31.00 ;
            RECT 129.00 24.00 131.00 26.00 ;
            RECT 129.00 19.00 131.00 21.00 ;
        END
    END selrom
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 138.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 79.00 29.00 125.00 31.00 ;
        RECT 79.00 69.00 125.00 71.00 ;
        RECT 4.00 74.00 136.00 76.00 ;
        RECT 4.00 24.00 136.00 26.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 44.00 19.00 51.00 21.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 44.00 79.00 51.00 81.00 ;
        RECT 64.00 19.00 96.00 21.00 ;
        RECT 64.00 79.00 96.00 81.00 ;
        RECT 4.00 79.00 136.00 81.00 ;
        RECT 4.00 19.00 136.00 21.00 ;
        RECT 119.00 74.00 136.00 76.00 ;
        RECT 119.00 24.00 136.00 26.00 ;
        RECT 9.00 39.00 45.00 41.00 ;
        RECT 4.00 39.00 46.00 41.00 ;
        RECT 4.00 59.00 26.00 61.00 ;
        RECT 9.00 59.00 26.00 61.00 ;
        RECT 59.00 24.00 81.00 26.00 ;
        RECT 19.00 24.00 41.00 26.00 ;
        RECT 19.00 74.00 41.00 76.00 ;
        RECT 59.00 74.00 81.00 76.00 ;
        RECT 4.00 69.00 136.00 71.00 ;
        RECT 4.00 29.00 136.00 31.00 ;
    END
END rom_dec_selmux23_ts


MACRO rom_dec_selmux45
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      120.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
            RECT 84.00 9.00 86.00 11.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
            RECT 74.00 9.00 76.00 11.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
            RECT 64.00 9.00 66.00 11.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 89.00 111.00 91.00 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 84.00 89.00 86.00 91.00 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 4.00 89.00 6.00 91.00 ;
            LAYER L_ALU3 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 104.00 84.00 106.00 86.00 ;
            RECT 104.00 79.00 106.00 81.00 ;
            RECT 104.00 74.00 106.00 76.00 ;
            RECT 104.00 69.00 106.00 71.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 104.00 59.00 106.00 61.00 ;
            RECT 104.00 54.00 106.00 56.00 ;
            RECT 104.00 49.00 106.00 51.00 ;
            RECT 104.00 44.00 106.00 46.00 ;
            RECT 104.00 39.00 106.00 41.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 104.00 29.00 106.00 31.00 ;
            RECT 104.00 24.00 106.00 26.00 ;
            RECT 104.00 19.00 106.00 21.00 ;
            RECT 104.00 14.00 106.00 16.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
        END
    END nck
    PIN sel4
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel4
    PIN sel5
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel5
    PIN mux4
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 74.00 39.00 76.00 41.00 ;
        END
    END mux4
    PIN mux5
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 54.00 59.00 56.00 61.00 ;
        END
    END mux5
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
            RECT 99.00 54.00 101.00 56.00 ;
            RECT 99.00 49.00 101.00 51.00 ;
            RECT 99.00 44.00 101.00 46.00 ;
            RECT 99.00 39.00 101.00 41.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
            RECT 99.00 14.00 101.00 16.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
        END
    END a5
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END selrom
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 74.00 116.00 76.00 ;
            RECT 114.00 69.00 116.00 71.00 ;
            RECT 114.00 64.00 116.00 66.00 ;
            RECT 114.00 59.00 116.00 61.00 ;
            RECT 114.00 54.00 116.00 56.00 ;
            RECT 114.00 49.00 116.00 51.00 ;
            RECT 114.00 44.00 116.00 46.00 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
        END
    END ck
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 118.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 39.00 79.00 46.00 81.00 ;
        RECT 39.00 19.00 46.00 21.00 ;
        RECT 9.00 59.00 56.00 61.00 ;
        RECT 9.00 39.00 75.00 41.00 ;
        RECT 79.00 69.00 111.00 71.00 ;
        RECT 29.00 74.00 41.00 76.00 ;
        RECT 59.00 74.00 91.00 76.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 59.00 24.00 91.00 26.00 ;
        RECT 29.00 24.00 41.00 26.00 ;
        RECT 79.00 29.00 111.00 31.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 64.00 19.00 101.00 21.00 ;
        RECT 64.00 79.00 101.00 81.00 ;
        RECT 4.00 19.00 116.00 21.00 ;
        RECT 4.00 24.00 116.00 26.00 ;
        RECT 4.00 29.00 116.00 31.00 ;
        RECT 4.00 39.00 116.00 41.00 ;
        RECT 4.00 59.00 116.00 61.00 ;
        RECT 4.00 69.00 116.00 71.00 ;
        RECT 4.00 74.00 116.00 76.00 ;
        RECT 4.00 79.00 116.00 81.00 ;
    END
END rom_dec_selmux45


MACRO rom_dec_selmux45_ts
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      140.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 109.00 89.00 111.00 91.00 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 84.00 89.00 86.00 91.00 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 4.00 89.00 6.00 91.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
            RECT 84.00 9.00 86.00 11.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
            RECT 74.00 9.00 76.00 11.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
            RECT 64.00 9.00 66.00 11.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
            LAYER L_ALU3 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 104.00 84.00 106.00 86.00 ;
            RECT 104.00 79.00 106.00 81.00 ;
            RECT 104.00 74.00 106.00 76.00 ;
            RECT 104.00 69.00 106.00 71.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 104.00 59.00 106.00 61.00 ;
            RECT 104.00 54.00 106.00 56.00 ;
            RECT 104.00 49.00 106.00 51.00 ;
            RECT 104.00 44.00 106.00 46.00 ;
            RECT 104.00 39.00 106.00 41.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 104.00 29.00 106.00 31.00 ;
            RECT 104.00 24.00 106.00 26.00 ;
            RECT 104.00 19.00 106.00 21.00 ;
            RECT 104.00 14.00 106.00 16.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
        END
    END nck
    PIN sel4
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel4
    PIN sel5
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel5
    PIN mux4
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 74.00 39.00 76.00 41.00 ;
        END
    END mux4
    PIN mux5
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 54.00 59.00 56.00 61.00 ;
        END
    END mux5
    PIN nenx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 119.00 74.00 121.00 76.00 ;
            RECT 119.00 69.00 121.00 71.00 ;
            RECT 119.00 64.00 121.00 66.00 ;
            RECT 119.00 59.00 121.00 61.00 ;
            RECT 119.00 54.00 121.00 56.00 ;
            RECT 119.00 49.00 121.00 51.00 ;
            RECT 119.00 44.00 121.00 46.00 ;
            RECT 119.00 39.00 121.00 41.00 ;
            RECT 119.00 34.00 121.00 36.00 ;
            RECT 119.00 29.00 121.00 31.00 ;
            RECT 119.00 24.00 121.00 26.00 ;
        END
    END nenx
    PIN enx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END enx
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
            RECT 99.00 54.00 101.00 56.00 ;
            RECT 99.00 49.00 101.00 51.00 ;
            RECT 99.00 44.00 101.00 46.00 ;
            RECT 99.00 39.00 101.00 41.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
        END
    END a5
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 129.00 79.00 131.00 81.00 ;
            RECT 129.00 74.00 131.00 76.00 ;
            RECT 129.00 69.00 131.00 71.00 ;
            RECT 129.00 64.00 131.00 66.00 ;
            RECT 129.00 59.00 131.00 61.00 ;
            RECT 129.00 54.00 131.00 56.00 ;
            RECT 129.00 49.00 131.00 51.00 ;
            RECT 129.00 44.00 131.00 46.00 ;
            RECT 129.00 39.00 131.00 41.00 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 129.00 29.00 131.00 31.00 ;
            RECT 129.00 24.00 131.00 26.00 ;
            RECT 129.00 19.00 131.00 21.00 ;
        END
    END selrom
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 74.00 116.00 76.00 ;
            RECT 114.00 69.00 116.00 71.00 ;
            RECT 114.00 64.00 116.00 66.00 ;
            RECT 114.00 59.00 116.00 61.00 ;
            RECT 114.00 54.00 116.00 56.00 ;
            RECT 114.00 49.00 116.00 51.00 ;
            RECT 114.00 44.00 116.00 46.00 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 138.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 69.00 136.00 71.00 ;
        RECT 4.00 29.00 136.00 31.00 ;
        RECT 79.00 29.00 125.00 31.00 ;
        RECT 79.00 69.00 125.00 71.00 ;
        RECT 64.00 79.00 101.00 81.00 ;
        RECT 64.00 19.00 101.00 21.00 ;
        RECT 39.00 79.00 46.00 81.00 ;
        RECT 39.00 19.00 46.00 21.00 ;
        RECT 4.00 39.00 76.00 41.00 ;
        RECT 9.00 39.00 76.00 41.00 ;
        RECT 4.00 59.00 56.00 61.00 ;
        RECT 9.00 59.00 56.00 61.00 ;
        RECT 4.00 74.00 136.00 76.00 ;
        RECT 4.00 24.00 136.00 26.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 29.00 24.00 41.00 26.00 ;
        RECT 59.00 24.00 91.00 26.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 59.00 74.00 91.00 76.00 ;
        RECT 29.00 74.00 41.00 76.00 ;
        RECT 4.00 79.00 136.00 81.00 ;
        RECT 4.00 19.00 136.00 21.00 ;
        RECT 119.00 74.00 136.00 76.00 ;
        RECT 119.00 24.00 136.00 26.00 ;
    END
END rom_dec_selmux45_ts


MACRO rom_dec_selmux67
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      120.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN mux6
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 39.00 36.00 41.00 ;
        END
    END mux6
    PIN mux7
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 59.00 16.00 61.00 ;
        END
    END mux7
    PIN sel7
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel7
    PIN sel6
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel6
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 104.00 84.00 106.00 86.00 ;
            RECT 104.00 79.00 106.00 81.00 ;
            RECT 104.00 74.00 106.00 76.00 ;
            RECT 104.00 69.00 106.00 71.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 104.00 59.00 106.00 61.00 ;
            RECT 104.00 54.00 106.00 56.00 ;
            RECT 104.00 49.00 106.00 51.00 ;
            RECT 104.00 44.00 106.00 46.00 ;
            RECT 104.00 39.00 106.00 41.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 104.00 29.00 106.00 31.00 ;
            RECT 104.00 24.00 106.00 26.00 ;
            RECT 104.00 19.00 106.00 21.00 ;
            RECT 104.00 14.00 106.00 16.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 89.00 111.00 91.00 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 84.00 89.00 86.00 91.00 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 4.00 89.00 6.00 91.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
            RECT 84.00 9.00 86.00 11.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
            RECT 74.00 9.00 76.00 11.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
            RECT 64.00 9.00 66.00 11.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END nck
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END selrom
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 74.00 116.00 76.00 ;
            RECT 114.00 69.00 116.00 71.00 ;
            RECT 114.00 64.00 116.00 66.00 ;
            RECT 114.00 59.00 116.00 61.00 ;
            RECT 114.00 54.00 116.00 56.00 ;
            RECT 114.00 49.00 116.00 51.00 ;
            RECT 114.00 44.00 116.00 46.00 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
        END
    END ck
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
            RECT 99.00 54.00 101.00 56.00 ;
            RECT 99.00 49.00 101.00 51.00 ;
            RECT 99.00 44.00 101.00 46.00 ;
            RECT 99.00 39.00 101.00 41.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
            RECT 99.00 14.00 101.00 16.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
        END
    END a5
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 118.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 79.00 116.00 81.00 ;
        RECT 4.00 74.00 116.00 76.00 ;
        RECT 4.00 69.00 116.00 71.00 ;
        RECT 4.00 59.00 116.00 61.00 ;
        RECT 4.00 39.00 116.00 41.00 ;
        RECT 4.00 29.00 116.00 31.00 ;
        RECT 4.00 24.00 116.00 26.00 ;
        RECT 4.00 19.00 116.00 21.00 ;
        RECT 64.00 79.00 101.00 81.00 ;
        RECT 64.00 19.00 100.00 21.00 ;
        RECT 39.00 79.00 46.00 81.00 ;
        RECT 39.00 19.00 46.00 21.00 ;
        RECT 79.00 69.00 111.00 71.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 79.00 29.00 111.00 31.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 9.00 59.00 24.00 61.00 ;
        RECT 9.00 39.00 35.00 41.00 ;
        RECT 59.00 24.00 81.00 26.00 ;
        RECT 59.00 74.00 81.00 76.00 ;
        RECT 19.00 74.00 41.00 76.00 ;
        RECT 19.00 24.00 41.00 26.00 ;
    END
END rom_dec_selmux67


MACRO rom_dec_selmux67_128
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      120.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN a6x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 84.00 64.00 86.00 66.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 74.00 64.00 76.00 66.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 64.00 64.00 66.00 66.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 54.00 64.00 56.00 66.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 44.00 64.00 46.00 66.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 34.00 64.00 36.00 66.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 24.00 64.00 26.00 66.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 14.00 64.00 16.00 66.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
        END
    END a6x
    PIN na6x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 84.00 34.00 86.00 36.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 74.00 34.00 76.00 36.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 64.00 34.00 66.00 36.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
        END
    END na6x
    PIN mux6
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 39.00 36.00 41.00 ;
        END
    END mux6
    PIN mux7
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 59.00 16.00 61.00 ;
        END
    END mux7
    PIN sel7
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel7
    PIN sel6
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel6
    PIN a6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
            RECT 114.00 19.00 116.00 21.00 ;
            RECT 114.00 14.00 116.00 16.00 ;
            RECT 114.00 9.00 116.00 11.00 ;
        END
    END a6
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END selrom
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
            RECT 99.00 54.00 101.00 56.00 ;
            RECT 99.00 49.00 101.00 51.00 ;
            RECT 99.00 44.00 101.00 46.00 ;
            RECT 99.00 39.00 101.00 41.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
            RECT 99.00 14.00 101.00 16.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
        END
    END a5
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 118.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 74.00 116.00 76.00 ;
        RECT 4.00 69.00 116.00 71.00 ;
        RECT 64.00 79.00 101.00 81.00 ;
        RECT 64.00 19.00 100.00 21.00 ;
        RECT 39.00 79.00 46.00 81.00 ;
        RECT 39.00 19.00 46.00 21.00 ;
        RECT 79.00 69.00 111.00 71.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 79.00 29.00 111.00 31.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 9.00 59.00 24.00 61.00 ;
        RECT 9.00 39.00 35.00 41.00 ;
        RECT 59.00 24.00 81.00 26.00 ;
        RECT 59.00 74.00 81.00 76.00 ;
        RECT 19.00 74.00 41.00 76.00 ;
        RECT 19.00 24.00 41.00 26.00 ;
        RECT 4.00 19.00 101.00 21.00 ;
        RECT 4.00 24.00 81.00 26.00 ;
        RECT 4.00 29.00 111.00 31.00 ;
        RECT 4.00 39.00 36.00 41.00 ;
        RECT 4.00 59.00 26.00 61.00 ;
        RECT 4.00 79.00 101.00 81.00 ;
        LAYER L_ALU3 ;
        RECT 114.00 34.00 116.00 76.00 ;
        RECT 114.00 34.00 116.00 76.00 ;
    END
END rom_dec_selmux67_128


MACRO rom_dec_selmux67_128_ts
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      140.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN a6x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 84.00 34.00 86.00 36.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 74.00 34.00 76.00 36.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 64.00 34.00 66.00 36.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
        END
    END a6x
    PIN na6x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 114.00 64.00 116.00 66.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 84.00 64.00 86.00 66.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 74.00 64.00 76.00 66.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 64.00 64.00 66.00 66.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 54.00 64.00 56.00 66.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 44.00 64.00 46.00 66.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 34.00 64.00 36.00 66.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 24.00 64.00 26.00 66.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 14.00 64.00 16.00 66.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
        END
    END na6x
    PIN mux6
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 39.00 36.00 41.00 ;
        END
    END mux6
    PIN mux7
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 59.00 16.00 61.00 ;
        END
    END mux7
    PIN sel7
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel7
    PIN sel6
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel6
    PIN nenx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 119.00 74.00 121.00 76.00 ;
            RECT 119.00 69.00 121.00 71.00 ;
            RECT 119.00 64.00 121.00 66.00 ;
            RECT 119.00 59.00 121.00 61.00 ;
            RECT 119.00 54.00 121.00 56.00 ;
            RECT 119.00 49.00 121.00 51.00 ;
            RECT 119.00 44.00 121.00 46.00 ;
            RECT 119.00 39.00 121.00 41.00 ;
            RECT 119.00 34.00 121.00 36.00 ;
            RECT 119.00 29.00 121.00 31.00 ;
            RECT 119.00 24.00 121.00 26.00 ;
        END
    END nenx
    PIN enx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END enx
    PIN a6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 94.00 116.00 96.00 ;
            RECT 114.00 89.00 116.00 91.00 ;
            RECT 114.00 84.00 116.00 86.00 ;
            RECT 114.00 79.00 116.00 81.00 ;
            RECT 114.00 74.00 116.00 76.00 ;
            RECT 114.00 69.00 116.00 71.00 ;
        END
    END a6
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
            RECT 99.00 54.00 101.00 56.00 ;
            RECT 99.00 49.00 101.00 51.00 ;
            RECT 99.00 44.00 101.00 46.00 ;
            RECT 99.00 39.00 101.00 41.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
            RECT 99.00 14.00 101.00 16.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
        END
    END a5
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 129.00 79.00 131.00 81.00 ;
            RECT 129.00 74.00 131.00 76.00 ;
            RECT 129.00 69.00 131.00 71.00 ;
            RECT 129.00 64.00 131.00 66.00 ;
            RECT 129.00 59.00 131.00 61.00 ;
            RECT 129.00 54.00 131.00 56.00 ;
            RECT 129.00 49.00 131.00 51.00 ;
            RECT 129.00 44.00 131.00 46.00 ;
            RECT 129.00 39.00 131.00 41.00 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 129.00 29.00 131.00 31.00 ;
            RECT 129.00 24.00 131.00 26.00 ;
            RECT 129.00 19.00 131.00 21.00 ;
        END
    END selrom
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 138.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 79.00 69.00 125.00 71.00 ;
        RECT 79.00 29.00 125.00 31.00 ;
        RECT 119.00 24.00 136.00 26.00 ;
        RECT 119.00 74.00 136.00 76.00 ;
        RECT 4.00 19.00 136.00 21.00 ;
        RECT 4.00 79.00 136.00 81.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 4.00 24.00 136.00 26.00 ;
        RECT 4.00 74.00 136.00 76.00 ;
        RECT 39.00 19.00 46.00 21.00 ;
        RECT 39.00 79.00 46.00 81.00 ;
        RECT 64.00 19.00 101.00 21.00 ;
        RECT 64.00 79.00 101.00 81.00 ;
        RECT 4.00 59.00 26.00 61.00 ;
        RECT 9.00 59.00 24.00 61.00 ;
        RECT 4.00 39.00 36.00 41.00 ;
        RECT 9.00 39.00 36.00 41.00 ;
        RECT 19.00 24.00 41.00 26.00 ;
        RECT 19.00 74.00 41.00 76.00 ;
        RECT 59.00 24.00 81.00 26.00 ;
        RECT 59.00 74.00 81.00 76.00 ;
        RECT 4.00 69.00 136.00 71.00 ;
        RECT 4.00 29.00 136.00 31.00 ;
        LAYER L_ALU3 ;
        RECT 114.00 24.00 116.00 66.00 ;
        RECT 114.00 24.00 116.00 66.00 ;
    END
END rom_dec_selmux67_128_ts


MACRO rom_dec_selmux67_ts
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      140.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN enx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 69.00 111.00 71.00 ;
            RECT 109.00 64.00 111.00 66.00 ;
            RECT 109.00 59.00 111.00 61.00 ;
            RECT 109.00 54.00 111.00 56.00 ;
            RECT 109.00 49.00 111.00 51.00 ;
            RECT 109.00 44.00 111.00 46.00 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
        END
    END enx
    PIN nenx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 119.00 74.00 121.00 76.00 ;
            RECT 119.00 69.00 121.00 71.00 ;
            RECT 119.00 64.00 121.00 66.00 ;
            RECT 119.00 59.00 121.00 61.00 ;
            RECT 119.00 54.00 121.00 56.00 ;
            RECT 119.00 49.00 121.00 51.00 ;
            RECT 119.00 44.00 121.00 46.00 ;
            RECT 119.00 39.00 121.00 41.00 ;
            RECT 119.00 34.00 121.00 36.00 ;
            RECT 119.00 29.00 121.00 31.00 ;
            RECT 119.00 24.00 121.00 26.00 ;
        END
    END nenx
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 109.00 89.00 111.00 91.00 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 84.00 89.00 86.00 91.00 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 4.00 89.00 6.00 91.00 ;
            LAYER L_ALU2 ;
            RECT 109.00 9.00 111.00 11.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
            RECT 84.00 9.00 86.00 11.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
            RECT 74.00 9.00 76.00 11.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
            RECT 64.00 9.00 66.00 11.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
            LAYER L_ALU3 ;
            RECT 104.00 89.00 106.00 91.00 ;
            RECT 104.00 84.00 106.00 86.00 ;
            RECT 104.00 79.00 106.00 81.00 ;
            RECT 104.00 74.00 106.00 76.00 ;
            RECT 104.00 69.00 106.00 71.00 ;
            RECT 104.00 64.00 106.00 66.00 ;
            RECT 104.00 59.00 106.00 61.00 ;
            RECT 104.00 54.00 106.00 56.00 ;
            RECT 104.00 49.00 106.00 51.00 ;
            RECT 104.00 44.00 106.00 46.00 ;
            RECT 104.00 39.00 106.00 41.00 ;
            RECT 104.00 34.00 106.00 36.00 ;
            RECT 104.00 29.00 106.00 31.00 ;
            RECT 104.00 24.00 106.00 26.00 ;
            RECT 104.00 19.00 106.00 21.00 ;
            RECT 104.00 14.00 106.00 16.00 ;
            RECT 104.00 9.00 106.00 11.00 ;
        END
    END nck
    PIN sel6
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END sel6
    PIN sel7
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 84.00 84.00 86.00 86.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 74.00 84.00 76.00 86.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 64.00 84.00 66.00 86.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 54.00 84.00 56.00 86.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 44.00 84.00 46.00 86.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
        END
    END sel7
    PIN mux7
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 59.00 16.00 61.00 ;
        END
    END mux7
    PIN mux6
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 39.00 36.00 41.00 ;
        END
    END mux6
    PIN selrom
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 129.00 79.00 131.00 81.00 ;
            RECT 129.00 74.00 131.00 76.00 ;
            RECT 129.00 69.00 131.00 71.00 ;
            RECT 129.00 64.00 131.00 66.00 ;
            RECT 129.00 59.00 131.00 61.00 ;
            RECT 129.00 54.00 131.00 56.00 ;
            RECT 129.00 49.00 131.00 51.00 ;
            RECT 129.00 44.00 131.00 46.00 ;
            RECT 129.00 39.00 131.00 41.00 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 129.00 29.00 131.00 31.00 ;
            RECT 129.00 24.00 131.00 26.00 ;
            RECT 129.00 19.00 131.00 21.00 ;
        END
    END selrom
    PIN a5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
            RECT 99.00 54.00 101.00 56.00 ;
            RECT 99.00 49.00 101.00 51.00 ;
            RECT 99.00 44.00 101.00 46.00 ;
            RECT 99.00 39.00 101.00 41.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
            RECT 99.00 14.00 101.00 16.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
        END
    END a5
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 79.00 84.00 81.00 86.00 ;
            RECT 79.00 79.00 81.00 81.00 ;
            RECT 79.00 74.00 81.00 76.00 ;
            RECT 79.00 69.00 81.00 71.00 ;
            RECT 79.00 64.00 81.00 66.00 ;
            RECT 79.00 59.00 81.00 61.00 ;
            RECT 79.00 54.00 81.00 56.00 ;
            RECT 79.00 49.00 81.00 51.00 ;
            RECT 79.00 44.00 81.00 46.00 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END a4
    PIN na4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 89.00 91.00 91.00 ;
            RECT 89.00 84.00 91.00 86.00 ;
            RECT 89.00 79.00 91.00 81.00 ;
            RECT 89.00 74.00 91.00 76.00 ;
            RECT 89.00 69.00 91.00 71.00 ;
            RECT 89.00 64.00 91.00 66.00 ;
            RECT 89.00 59.00 91.00 61.00 ;
            RECT 89.00 54.00 91.00 56.00 ;
            RECT 89.00 49.00 91.00 51.00 ;
            RECT 89.00 44.00 91.00 46.00 ;
            RECT 89.00 39.00 91.00 41.00 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
            RECT 89.00 9.00 91.00 11.00 ;
        END
    END na4
    PIN na3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 69.00 84.00 71.00 86.00 ;
            RECT 69.00 79.00 71.00 81.00 ;
            RECT 69.00 74.00 71.00 76.00 ;
            RECT 69.00 69.00 71.00 71.00 ;
            RECT 69.00 64.00 71.00 66.00 ;
            RECT 69.00 59.00 71.00 61.00 ;
            RECT 69.00 54.00 71.00 56.00 ;
            RECT 69.00 49.00 71.00 51.00 ;
            RECT 69.00 44.00 71.00 46.00 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END na3
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 59.00 84.00 61.00 86.00 ;
            RECT 59.00 79.00 61.00 81.00 ;
            RECT 59.00 74.00 61.00 76.00 ;
            RECT 59.00 69.00 61.00 71.00 ;
            RECT 59.00 64.00 61.00 66.00 ;
            RECT 59.00 59.00 61.00 61.00 ;
            RECT 59.00 54.00 61.00 56.00 ;
            RECT 59.00 49.00 61.00 51.00 ;
            RECT 59.00 44.00 61.00 46.00 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END a3
    PIN na2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 49.00 84.00 51.00 86.00 ;
            RECT 49.00 79.00 51.00 81.00 ;
            RECT 49.00 74.00 51.00 76.00 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END na2
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 39.00 84.00 41.00 86.00 ;
            RECT 39.00 79.00 41.00 81.00 ;
            RECT 39.00 74.00 41.00 76.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 39.00 64.00 41.00 66.00 ;
            RECT 39.00 59.00 41.00 61.00 ;
            RECT 39.00 54.00 41.00 56.00 ;
            RECT 39.00 49.00 41.00 51.00 ;
            RECT 39.00 44.00 41.00 46.00 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END a2
    PIN na1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 29.00 84.00 31.00 86.00 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END na1
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
            RECT 19.00 64.00 21.00 66.00 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END a1
    PIN na0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END na0
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a0
    PIN na5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 89.00 96.00 91.00 ;
            RECT 94.00 84.00 96.00 86.00 ;
            RECT 94.00 79.00 96.00 81.00 ;
            RECT 94.00 74.00 96.00 76.00 ;
            RECT 94.00 69.00 96.00 71.00 ;
            RECT 94.00 64.00 96.00 66.00 ;
            RECT 94.00 59.00 96.00 61.00 ;
            RECT 94.00 54.00 96.00 56.00 ;
            RECT 94.00 49.00 96.00 51.00 ;
            RECT 94.00 44.00 96.00 46.00 ;
            RECT 94.00 39.00 96.00 41.00 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
            RECT 94.00 9.00 96.00 11.00 ;
        END
    END na5
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 74.00 116.00 76.00 ;
            RECT 114.00 69.00 116.00 71.00 ;
            RECT 114.00 64.00 116.00 66.00 ;
            RECT 114.00 59.00 116.00 61.00 ;
            RECT 114.00 54.00 116.00 56.00 ;
            RECT 114.00 49.00 116.00 51.00 ;
            RECT 114.00 44.00 116.00 46.00 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
        END
    END ck
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
    END vdd
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 1.50 138.50 98.50 ;
        LAYER L_ALU2 ;
        RECT 4.00 29.00 136.00 31.00 ;
        RECT 4.00 69.00 136.00 71.00 ;
        RECT 59.00 74.00 81.00 76.00 ;
        RECT 59.00 24.00 81.00 26.00 ;
        RECT 19.00 74.00 41.00 76.00 ;
        RECT 19.00 24.00 41.00 26.00 ;
        RECT 9.00 39.00 36.00 41.00 ;
        RECT 4.00 39.00 36.00 41.00 ;
        RECT 9.00 59.00 24.00 61.00 ;
        RECT 4.00 59.00 26.00 61.00 ;
        RECT 64.00 79.00 101.00 81.00 ;
        RECT 64.00 19.00 101.00 21.00 ;
        RECT 39.00 79.00 46.00 81.00 ;
        RECT 39.00 19.00 46.00 21.00 ;
        RECT 4.00 74.00 136.00 76.00 ;
        RECT 4.00 24.00 136.00 26.00 ;
        RECT 54.00 29.00 71.00 31.00 ;
        RECT 9.00 29.00 36.00 31.00 ;
        RECT 54.00 69.00 61.00 71.00 ;
        RECT 4.00 69.00 36.00 71.00 ;
        RECT 4.00 79.00 136.00 81.00 ;
        RECT 4.00 19.00 136.00 21.00 ;
        RECT 119.00 74.00 136.00 76.00 ;
        RECT 119.00 24.00 136.00 26.00 ;
        RECT 79.00 29.00 125.00 31.00 ;
        RECT 79.00 69.00 125.00 71.00 ;
    END
END rom_dec_selmux67_ts


END LIBRARY
