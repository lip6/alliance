#
# $Id: cmos.lef,v 1.2 2002/10/03 17:14:02 xtof Exp $
#
# /------------------------------------------------------------------\
# |                                                                  |
# |        A l l i a n c e   C A D   S y s t e m                     |
# |  S i l i c o n   E n s e m b l e / A l l i a n c e               |
# |                                                                  |
# |  Author    :                      Jean-Paul CHAPUT               |
# |  E-mail    :         alliance-users@asim.lip6.fr               |
# | ================================================================ |
# |  LEF       :         "./cmos_12.lef"                             |
# | **************************************************************** |
# |  U p d a t e s                                                   |
# |                                                                  |
# \------------------------------------------------------------------/
#

VERSION 5.1 ;

NAMESCASESENSITIVE    ON ;

#NOWIREEXTENSIONATPIN ON ;


UNITS
    DATABASE MICRONS 100  ;
END UNITS


LAYER L_POLY
    TYPE MASTERSLICE ;
END L_POLY


LAYER L_CONT
    TYPE CUT ;
END L_CONT


LAYER L_ALU1
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END L_ALU1


LAYER L_VIA1
    TYPE CUT ;
END L_VIA1


LAYER L_ALU2
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END L_ALU2


LAYER L_VIA2
    TYPE CUT ;
END L_VIA2


LAYER L_ALU3
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END L_ALU3


LAYER L_VIA3
    TYPE CUT ;
END L_VIA3


LAYER L_ALU4
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END L_ALU4


LAYER L_VIA4
    TYPE CUT ;
END L_VIA4


LAYER L_ALU5
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END L_ALU5


LAYER L_VIA5
    TYPE CUT ;
END L_VIA5


LAYER L_ALU6
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END L_ALU6


#VIA CONT_POLY DEFAULT
#    LAYER L_POLY ;
#        RECT -1.50 -1.50 1.50 1.50 ;
#    LAYER L_CONT ;
#        RECT -0.50 -0.50 0.50 0.50 ;
#    LAYER L_ALU1 ;
#        RECT -1.00 -1.00 1.00 1.00 ;
#END CONT_POLY


VIA CONT_VIA DEFAULT
    LAYER L_ALU1 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER L_VIA1 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER L_ALU2 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA


VIA CONT_VIA2 DEFAULT
    LAYER L_ALU3 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER L_VIA2 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER L_ALU2 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA2


VIA CONT_VIA3 DEFAULT
    LAYER L_ALU4 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER L_VIA3 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER L_ALU3 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA3


VIA CONT_VIA4 DEFAULT
    LAYER L_ALU5 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER L_VIA4 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER L_ALU4 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA4


VIA CONT_VIA5 DEFAULT
    LAYER L_ALU6 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER L_VIA5 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER L_ALU5 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA5


VIARULE TURN_ALU1 GENERATE
    LAYER L_ALU1 ;
        DIRECTION vertical ;

    LAYER L_ALU1 ;
        DIRECTION horizontal ;
END TURN_ALU1


VIARULE TURN_ALU2 GENERATE
    LAYER L_ALU2 ;
        DIRECTION vertical ;

    LAYER L_ALU2 ;
        DIRECTION horizontal ;
END TURN_ALU2


VIARULE TURN_ALU3 GENERATE
    LAYER L_ALU3 ;
        DIRECTION vertical ;

    LAYER L_ALU3 ;
        DIRECTION horizontal ;
END TURN_ALU3


VIARULE TURN_ALU4 GENERATE
    LAYER L_ALU4 ;
        DIRECTION vertical ;

    LAYER L_ALU4 ;
        DIRECTION horizontal ;
END TURN_ALU4


VIARULE TURN_ALU5 GENERATE
    LAYER L_ALU5 ;
        DIRECTION vertical ;

    LAYER L_ALU5 ;
        DIRECTION horizontal ;
END TURN_ALU5


VIARULE TURN_ALU6 GENERATE
    LAYER L_ALU6 ;
        DIRECTION vertical ;

    LAYER L_ALU6 ;
        DIRECTION horizontal ;
END TURN_ALU6


#VIARULE VIA1_HV
#    LAYER L_ALU1 ;
#        DIRECTION VERTICAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    LAYER L_ALU2 ;
#        DIRECTION HORIZONTAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    VIA CONT_VIA ;
#END VIA1_HV
#
#
#VIARULE VIA2_VH
#    LAYER L_ALU2 ;
#        DIRECTION HORIZONTAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    LAYER L_ALU3 ;
#        DIRECTION VERTICAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    VIA CONT_VIA2 ;
#END VIA2_VH
#
#
#VIARULE VIA3_VH
#    LAYER L_ALU3 ;
#        DIRECTION HORIZONTAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    LAYER L_ALU4 ;
#        DIRECTION VERTICAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    VIA CONT_VIA3 ;
#END VIA3_VH


VIARULE genVIA1_HV GENERATE
    LAYER L_ALU1 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_ALU2 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_VIA1 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA1_HV


VIARULE genVIA1_VH GENERATE
    LAYER L_ALU1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_ALU2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_VIA1 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA1_VH


VIARULE genVIA2_VH GENERATE
    LAYER L_ALU2 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_ALU3 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_VIA2 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA2_VH


VIARULE genVIA2_HV GENERATE
    LAYER L_ALU2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_ALU3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_VIA2 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA2_HV


VIARULE genVIA3_VH GENERATE
    LAYER L_ALU3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_ALU4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_VIA3 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA3_VH


VIARULE genVIA3_HV GENERATE
    LAYER L_ALU3 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_ALU4 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER L_VIA3 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA3_HV


SPACING
    SAMENET L_CONT L_CONT 3.00 ;
    SAMENET L_VIA1 L_VIA1 3.00 ;
    SAMENET L_VIA2 L_VIA2 3.00 ;
    SAMENET L_CONT L_VIA1 3.00 STACK ;
    SAMENET L_VIA1 L_VIA2 3.00 STACK ;
    SAMENET L_VIA2 L_VIA3 3.00 STACK ;
    SAMENET L_VIA3 L_VIA4 3.00 STACK ;
    SAMENET L_VIA4 L_VIA5 3.00 STACK ;
    SAMENET L_POLY L_POLY 3.00 ;
    SAMENET L_ALU1 L_ALU1 3.00 STACK ;
    SAMENET L_ALU2 L_ALU2 3.00 STACK ;
    SAMENET L_ALU3 L_ALU3 3.00 STACK ;
    SAMENET L_ALU4 L_ALU4 3.00 STACK ;
    SAMENET L_ALU5 L_ALU5 3.00 STACK ;
    SAMENET L_ALU6 L_ALU6 3.00 ;
END SPACING


SITE core
    SYMMETRY y  ;
    CLASS core  ;
    SIZE 5.00 BY 50.00 ;
END core


SITE pad
    SYMMETRY y  ;
    CLASS pad  ;
    SIZE 1.00 BY 500.00 ;
END pad


SITE corner
    SYMMETRY y r90  ;
    CLASS pad  ;
    SIZE 500.00 BY 500.00 ;
END corner


END LIBRARY
