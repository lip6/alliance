
MACRO rf_dec_bufad0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END nq
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 29.00 26.00 31.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 10.00 6.00 10.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 43.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 43.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 43.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 43.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 43.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 43.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 43.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 -1.00 16.00 1.00 ;
    END
END rf_dec_bufad0


MACRO rf_dec_bufad1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END nq
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 10.00 6.00 10.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 31.00 21.00 ;
        RECT 4.00 -1.00 16.00 1.00 ;
    END
END rf_dec_bufad1


MACRO rf_dec_bufad1r
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END q
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 10.00 6.00 10.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 31.00 21.00 ;
        RECT 4.00 49.00 16.00 51.00 ;
    END
END rf_dec_bufad1r


MACRO rf_dec_bufad2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq1
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END nq1
    PIN nq0
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END nq0
    PIN q1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END q1
    PIN q0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END q0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 10.00 6.00 10.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 46.00 21.00 ;
        RECT 4.00 -1.00 16.00 1.00 ;
    END
END rf_dec_bufad2


MACRO rf_dec_bufad2r
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq1
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END nq1
    PIN nq0
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END nq0
    PIN q1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END q1
    PIN q0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END q0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 10.00 6.00 10.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 46.00 21.00 ;
        RECT 4.00 49.00 16.00 51.00 ;
    END
END rf_dec_bufad2r


MACRO rf_dec_nand2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 36.00 21.00 ;
    END
END rf_dec_nand2


MACRO rf_dec_nand3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 29.00 19.00 36.00 21.00 ;
        RECT 19.00 19.00 41.00 21.00 ;
    END
END rf_dec_nand3


MACRO rf_dec_nand4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END nq
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i0
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 14.00 19.00 41.00 21.00 ;
        RECT 29.00 19.00 36.00 21.00 ;
    END
END rf_dec_nand4


MACRO rf_dec_nao3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END nq
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 34.00 21.00 36.00 ;
        END
    END i2
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 39.00 11.00 41.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 23.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 23.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 23.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 23.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 23.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 23.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 23.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 19.00 11.00 21.00 ;
    END
END rf_dec_nao3


MACRO rf_dec_nbuf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      55.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 52.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 45.00 6.00 45.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 52.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 53.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 53.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 53.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 53.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 53.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 53.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 53.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 39.00 49.00 51.00 51.00 ;
    END
END rf_dec_nbuf


MACRO rf_dec_nor3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 39.00 11.00 41.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 23.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 23.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 23.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 23.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 23.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 23.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 23.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 19.00 11.00 21.00 ;
    END
END rf_dec_nor3


MACRO rf_fifo_buf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN nreset
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 59.00 46.00 61.00 ;
            RECT 44.00 54.00 46.00 56.00 ;
            RECT 44.00 49.00 46.00 51.00 ;
            RECT 44.00 44.00 46.00 46.00 ;
            RECT 44.00 39.00 46.00 41.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
        END
    END nreset
    PIN xreset
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END xreset
    PIN nr
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT 4.00 84.00 6.00 86.00 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
            RECT 4.00 59.00 6.00 61.00 ;
        END
    END nr
    PIN nw
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 24.00 79.00 26.00 81.00 ;
            RECT 24.00 74.00 26.00 76.00 ;
            RECT 24.00 69.00 26.00 71.00 ;
            RECT 24.00 64.00 26.00 66.00 ;
            RECT 24.00 59.00 26.00 61.00 ;
        END
    END nw
    PIN xckm
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 39.00 36.00 41.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
        END
    END xckm
    PIN xcks
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END xcks
    PIN reset
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 79.00 41.00 81.00 ;
        END
    END reset
    PIN cks
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 39.00 21.00 41.00 ;
        END
    END cks
    PIN ckm
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END ckm
    PIN r
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 84.00 11.00 86.00 ;
        END
    END r
    PIN w
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 74.00 31.00 76.00 ;
        END
    END w
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 47.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 47.00 97.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 21.00 61.00 ;
        RECT 24.00 59.00 26.00 61.00 ;
        RECT 29.00 59.00 31.00 61.00 ;
        RECT 34.00 59.00 36.00 61.00 ;
        RECT 39.00 59.00 41.00 61.00 ;
        RECT 44.00 59.00 48.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 26.00 66.00 ;
        RECT 29.00 64.00 31.00 66.00 ;
        RECT 34.00 64.00 36.00 66.00 ;
        RECT 39.00 64.00 41.00 66.00 ;
        RECT 44.00 64.00 48.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 21.00 71.00 ;
        RECT 24.00 69.00 26.00 71.00 ;
        RECT 29.00 69.00 31.00 71.00 ;
        RECT 34.00 69.00 36.00 71.00 ;
        RECT 39.00 69.00 41.00 71.00 ;
        RECT 44.00 69.00 48.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 21.00 76.00 ;
        RECT 24.00 74.00 26.00 76.00 ;
        RECT 29.00 74.00 31.00 76.00 ;
        RECT 34.00 74.00 36.00 76.00 ;
        RECT 39.00 74.00 41.00 76.00 ;
        RECT 44.00 74.00 48.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 21.00 81.00 ;
        RECT 24.00 79.00 26.00 81.00 ;
        RECT 29.00 79.00 31.00 81.00 ;
        RECT 34.00 79.00 36.00 81.00 ;
        RECT 39.00 79.00 41.00 81.00 ;
        RECT 44.00 79.00 48.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 21.00 86.00 ;
        RECT 24.00 84.00 26.00 86.00 ;
        RECT 29.00 84.00 31.00 86.00 ;
        RECT 34.00 84.00 36.00 86.00 ;
        RECT 39.00 84.00 41.00 86.00 ;
        RECT 44.00 84.00 48.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 21.00 91.00 ;
        RECT 24.00 89.00 26.00 91.00 ;
        RECT 29.00 89.00 31.00 91.00 ;
        RECT 34.00 89.00 36.00 91.00 ;
        RECT 39.00 89.00 41.00 91.00 ;
        RECT 44.00 89.00 48.50 91.00 ;
        LAYER L_ALU2 ;
        RECT 44.00 24.00 51.00 26.00 ;
        RECT 44.00 59.00 51.00 61.00 ;
    END
END rf_fifo_buf


MACRO rf_fifo_clock
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN ckm
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
            RECT 9.00 54.00 11.00 56.00 ;
            RECT 9.00 49.00 11.00 51.00 ;
            RECT 9.00 44.00 11.00 46.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
        END
    END ckm
    PIN cks
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 79.00 31.00 81.00 ;
            RECT 29.00 74.00 31.00 76.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 29.00 64.00 31.00 66.00 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
        END
    END cks
    PIN ckok
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 9.00 84.00 11.00 86.00 ;
            RECT 9.00 79.00 11.00 81.00 ;
            RECT 9.00 74.00 11.00 76.00 ;
            RECT 9.00 69.00 11.00 71.00 ;
            RECT 9.00 64.00 11.00 66.00 ;
            RECT 9.00 59.00 11.00 61.00 ;
        END
    END ckok
    PIN wok
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 79.00 6.00 81.00 ;
            RECT 4.00 74.00 6.00 76.00 ;
            RECT 4.00 69.00 6.00 71.00 ;
            RECT 4.00 64.00 6.00 66.00 ;
        END
    END wok
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 49.00 64.00 51.00 66.00 ;
            RECT 49.00 59.00 51.00 61.00 ;
            RECT 49.00 54.00 51.00 56.00 ;
            RECT 49.00 49.00 51.00 51.00 ;
            RECT 49.00 44.00 51.00 46.00 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            LAYER L_ALU2 ;
            RECT 49.00 69.00 51.00 71.00 ;
            RECT 44.00 69.00 46.00 71.00 ;
            RECT 39.00 69.00 41.00 71.00 ;
            RECT 34.00 69.00 36.00 71.00 ;
            RECT 29.00 69.00 31.00 71.00 ;
            RECT 24.00 69.00 26.00 71.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
        END
    END ck
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 47.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 47.00 97.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 21.00 61.00 ;
        RECT 24.00 59.00 26.00 61.00 ;
        RECT 29.00 59.00 31.00 61.00 ;
        RECT 34.00 59.00 36.00 61.00 ;
        RECT 39.00 59.00 41.00 61.00 ;
        RECT 44.00 59.00 48.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 26.00 66.00 ;
        RECT 29.00 64.00 31.00 66.00 ;
        RECT 34.00 64.00 36.00 66.00 ;
        RECT 39.00 64.00 41.00 66.00 ;
        RECT 44.00 64.00 48.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 21.00 71.00 ;
        RECT 24.00 69.00 26.00 71.00 ;
        RECT 29.00 69.00 31.00 71.00 ;
        RECT 34.00 69.00 36.00 71.00 ;
        RECT 39.00 69.00 41.00 71.00 ;
        RECT 44.00 69.00 48.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 21.00 76.00 ;
        RECT 24.00 74.00 26.00 76.00 ;
        RECT 29.00 74.00 31.00 76.00 ;
        RECT 34.00 74.00 36.00 76.00 ;
        RECT 39.00 74.00 41.00 76.00 ;
        RECT 44.00 74.00 48.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 21.00 81.00 ;
        RECT 24.00 79.00 26.00 81.00 ;
        RECT 29.00 79.00 31.00 81.00 ;
        RECT 34.00 79.00 36.00 81.00 ;
        RECT 39.00 79.00 41.00 81.00 ;
        RECT 44.00 79.00 48.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 21.00 86.00 ;
        RECT 24.00 84.00 26.00 86.00 ;
        RECT 29.00 84.00 31.00 86.00 ;
        RECT 34.00 84.00 36.00 86.00 ;
        RECT 39.00 84.00 41.00 86.00 ;
        RECT 44.00 84.00 48.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 21.00 91.00 ;
        RECT 24.00 89.00 26.00 91.00 ;
        RECT 29.00 89.00 31.00 91.00 ;
        RECT 34.00 89.00 36.00 91.00 ;
        RECT 39.00 89.00 41.00 91.00 ;
        RECT 44.00 89.00 48.50 91.00 ;
        LAYER L_ALU2 ;
        RECT 9.00 24.00 51.00 26.00 ;
        RECT 9.00 39.00 16.00 41.00 ;
        RECT 24.00 39.00 31.00 41.00 ;
        RECT 29.00 19.00 41.00 21.00 ;
        RECT 9.00 24.00 36.00 26.00 ;
        RECT 34.00 59.00 41.00 61.00 ;
        RECT 9.00 84.00 36.00 86.00 ;
        RECT 29.00 79.00 46.00 81.00 ;
        RECT 9.00 84.00 36.00 86.00 ;
        RECT 29.00 19.00 41.00 21.00 ;
        RECT 9.00 39.00 46.00 41.00 ;
        LAYER L_ALU3 ;
        RECT 39.00 19.00 41.00 61.00 ;
        RECT 34.00 24.00 36.00 61.00 ;
        RECT 44.00 39.00 46.00 81.00 ;
        RECT 44.00 39.00 46.00 81.00 ;
        RECT 34.00 24.00 36.00 61.00 ;
        RECT 39.00 19.00 41.00 61.00 ;
    END
END rf_fifo_clock


MACRO rf_fifo_empty
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN empty
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 39.00 46.00 41.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
        END
    END empty
    PIN emptynext
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 29.00 11.00 31.00 ;
        END
    END emptynext
    PIN nreset
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END nreset
    PIN ckm
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END ckm
    PIN cks
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END cks
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
    END
END rf_fifo_empty


MACRO rf_fifo_full
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN full
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 39.00 46.00 41.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
        END
    END full
    PIN reset
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END reset
    PIN ckm
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END ckm
    PIN cks
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END cks
    PIN fullnext
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 24.00 11.00 26.00 ;
        END
    END fullnext
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
    END
END rf_fifo_full


MACRO rf_fifo_inc
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN inc
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 4.00 39.00 6.00 41.00 ;
        END
    END inc
    PIN ckm
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END ckm
    PIN nreset
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 24.00 21.00 26.00 ;
        END
    END nreset
    PIN nval
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 39.00 31.00 41.00 ;
        END
    END nval
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
    END
END rf_fifo_inc


MACRO rf_fifo_nop
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nval
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 39.00 31.00 41.00 ;
        END
    END nval
    PIN nop
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 4.00 39.00 6.00 41.00 ;
        END
    END nop
    PIN rwok
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 29.00 41.00 31.00 ;
        END
    END rwok
    PIN rw
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 44.00 14.00 46.00 16.00 ;
        END
    END rw
    PIN nreset
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 24.00 21.00 26.00 ;
        END
    END nreset
    PIN ckm
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END ckm
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
    END
END rf_fifo_nop


MACRO rf_fifo_ok
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN ok
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END ok
    PIN nextval
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 29.00 16.00 31.00 ;
        END
    END nextval
    PIN ripple
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 44.00 34.00 46.00 36.00 ;
        END
    END ripple
    PIN nrw
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END nrw
    PIN rw
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 24.00 36.00 26.00 ;
        END
    END rw
    PIN prev
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END prev
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
    END
END rf_fifo_ok


MACRO rf_fifo_orand4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN rippleout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END rippleout
    PIN b1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END b1
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END a1
    PIN b0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END b0
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
        END
    END a0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
    END
END rf_fifo_orand4


MACRO rf_fifo_orand5
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN rippleout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END rippleout
    PIN b1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END b1
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END a1
    PIN b0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
        END
    END b0
    PIN a0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END a0
    PIN ripplein
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END ripplein
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
    END
END rf_fifo_orand5


MACRO rf_fifo_ptreset
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN pt
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END pt
    PIN cks
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END cks
    PIN nop
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END nop
    PIN reset
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END reset
    PIN inc
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END inc
    PIN ptm1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END ptm1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 34.00 41.00 36.00 ;
        RECT 4.00 34.00 41.00 36.00 ;
        RECT 34.00 19.00 41.00 21.00 ;
        RECT 9.00 19.00 16.00 21.00 ;
        RECT 9.00 19.00 41.00 21.00 ;
    END
END rf_fifo_ptreset


MACRO rf_fifo_ptset
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN pt
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 44.00 9.00 46.00 11.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END pt
    PIN nop
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END nop
    PIN ptm1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END ptm1
    PIN nreset
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END nreset
    PIN cks
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END cks
    PIN inc
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END inc
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 9.00 19.00 16.00 21.00 ;
        RECT 34.00 19.00 41.00 21.00 ;
        RECT 4.00 34.00 41.00 36.00 ;
        RECT 9.00 19.00 41.00 21.00 ;
        RECT 4.00 34.00 41.00 36.00 ;
    END
END rf_fifo_ptset


MACRO rf_inmux_buf_2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 89.00 36.00 91.00 ;
        END
    END nck
    PIN sel0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 39.00 36.00 41.00 ;
        END
    END sel0
    PIN sel1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END sel1
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
        END
    END ck
    PIN sel
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 14.00 79.00 16.00 81.00 ;
            RECT 14.00 74.00 16.00 76.00 ;
            RECT 14.00 69.00 16.00 71.00 ;
        END
    END sel
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 42.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 42.00 97.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 10.00 6.00 10.00 94.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 43.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 43.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 43.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 43.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 43.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 43.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 43.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 21.00 61.00 ;
        RECT 24.00 59.00 26.00 61.00 ;
        RECT 29.00 59.00 31.00 61.00 ;
        RECT 34.00 59.00 36.00 61.00 ;
        RECT 39.00 59.00 43.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 26.00 66.00 ;
        RECT 29.00 64.00 31.00 66.00 ;
        RECT 34.00 64.00 36.00 66.00 ;
        RECT 39.00 64.00 43.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 21.00 71.00 ;
        RECT 24.00 69.00 26.00 71.00 ;
        RECT 29.00 69.00 31.00 71.00 ;
        RECT 34.00 69.00 36.00 71.00 ;
        RECT 39.00 69.00 43.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 21.00 76.00 ;
        RECT 24.00 74.00 26.00 76.00 ;
        RECT 29.00 74.00 31.00 76.00 ;
        RECT 34.00 74.00 36.00 76.00 ;
        RECT 39.00 74.00 43.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 21.00 81.00 ;
        RECT 24.00 79.00 26.00 81.00 ;
        RECT 29.00 79.00 31.00 81.00 ;
        RECT 34.00 79.00 36.00 81.00 ;
        RECT 39.00 79.00 43.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 21.00 86.00 ;
        RECT 24.00 84.00 26.00 86.00 ;
        RECT 29.00 84.00 31.00 86.00 ;
        RECT 34.00 84.00 36.00 86.00 ;
        RECT 39.00 84.00 43.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 21.00 91.00 ;
        RECT 24.00 89.00 26.00 91.00 ;
        RECT 29.00 89.00 31.00 91.00 ;
        RECT 34.00 89.00 36.00 91.00 ;
        RECT 39.00 89.00 43.50 91.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 99.00 16.00 101.00 ;
        RECT 4.00 -1.00 16.00 1.00 ;
        RECT 26.00 39.00 40.00 41.00 ;
        RECT 8.00 14.00 26.00 16.00 ;
        RECT 4.00 14.00 26.00 16.00 ;
        RECT 24.00 39.00 41.00 41.00 ;
    END
END rf_inmux_buf_2


MACRO rf_inmux_buf_4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 200.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN sel1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 184.00 26.00 186.00 ;
            RECT 24.00 179.00 26.00 181.00 ;
            RECT 24.00 174.00 26.00 176.00 ;
            RECT 24.00 169.00 26.00 171.00 ;
            RECT 24.00 164.00 26.00 166.00 ;
            RECT 24.00 159.00 26.00 161.00 ;
            RECT 24.00 154.00 26.00 156.00 ;
            RECT 24.00 149.00 26.00 151.00 ;
            RECT 24.00 144.00 26.00 146.00 ;
            RECT 24.00 139.00 26.00 141.00 ;
            RECT 24.00 134.00 26.00 136.00 ;
            RECT 24.00 129.00 26.00 131.00 ;
            RECT 24.00 124.00 26.00 126.00 ;
            RECT 24.00 119.00 26.00 121.00 ;
            RECT 24.00 114.00 26.00 116.00 ;
            RECT 24.00 109.00 26.00 111.00 ;
            RECT 24.00 104.00 26.00 106.00 ;
            RECT 24.00 99.00 26.00 101.00 ;
            RECT 24.00 94.00 26.00 96.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 24.00 84.00 26.00 86.00 ;
            RECT 24.00 79.00 26.00 81.00 ;
            RECT 24.00 74.00 26.00 76.00 ;
            RECT 24.00 69.00 26.00 71.00 ;
            RECT 24.00 64.00 26.00 66.00 ;
            RECT 24.00 59.00 26.00 61.00 ;
            RECT 24.00 54.00 26.00 56.00 ;
            RECT 24.00 49.00 26.00 51.00 ;
            RECT 24.00 44.00 26.00 46.00 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END sel1
    PIN sel0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 159.00 36.00 161.00 ;
            RECT 34.00 154.00 36.00 156.00 ;
            RECT 34.00 149.00 36.00 151.00 ;
            RECT 34.00 144.00 36.00 146.00 ;
            RECT 34.00 139.00 36.00 141.00 ;
            RECT 34.00 134.00 36.00 136.00 ;
            RECT 34.00 129.00 36.00 131.00 ;
            RECT 34.00 124.00 36.00 126.00 ;
            RECT 34.00 119.00 36.00 121.00 ;
            RECT 34.00 114.00 36.00 116.00 ;
            RECT 34.00 109.00 36.00 111.00 ;
            RECT 34.00 104.00 36.00 106.00 ;
            RECT 34.00 99.00 36.00 101.00 ;
            RECT 34.00 94.00 36.00 96.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 34.00 84.00 36.00 86.00 ;
            RECT 34.00 79.00 36.00 81.00 ;
            RECT 34.00 74.00 36.00 76.00 ;
            RECT 34.00 69.00 36.00 71.00 ;
            RECT 34.00 64.00 36.00 66.00 ;
            RECT 34.00 59.00 36.00 61.00 ;
            RECT 34.00 54.00 36.00 56.00 ;
            RECT 34.00 49.00 36.00 51.00 ;
            RECT 34.00 44.00 36.00 46.00 ;
            RECT 34.00 39.00 36.00 41.00 ;
        END
    END sel0
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
        END
    END nck
    PIN sel
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 14.00 79.00 16.00 81.00 ;
            RECT 14.00 74.00 16.00 76.00 ;
            RECT 14.00 69.00 16.00 71.00 ;
        END
    END sel
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 19.00 84.00 21.00 86.00 ;
            RECT 19.00 79.00 21.00 81.00 ;
            RECT 19.00 74.00 21.00 76.00 ;
            RECT 19.00 69.00 21.00 71.00 ;
        END
    END ck
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 42.00 53.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 147.00 42.00 147.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 153.00 42.00 153.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 42.00 97.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 103.00 42.00 103.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 197.00 42.00 197.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 10.00 6.00 10.00 194.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 43.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 43.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 43.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 43.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 43.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 43.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 43.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 21.00 61.00 ;
        RECT 24.00 59.00 26.00 61.00 ;
        RECT 29.00 59.00 31.00 61.00 ;
        RECT 34.00 59.00 36.00 61.00 ;
        RECT 39.00 59.00 43.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 26.00 66.00 ;
        RECT 29.00 64.00 31.00 66.00 ;
        RECT 34.00 64.00 36.00 66.00 ;
        RECT 39.00 64.00 43.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 21.00 71.00 ;
        RECT 24.00 69.00 26.00 71.00 ;
        RECT 29.00 69.00 31.00 71.00 ;
        RECT 34.00 69.00 36.00 71.00 ;
        RECT 39.00 69.00 43.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 21.00 76.00 ;
        RECT 24.00 74.00 26.00 76.00 ;
        RECT 29.00 74.00 31.00 76.00 ;
        RECT 34.00 74.00 36.00 76.00 ;
        RECT 39.00 74.00 43.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 21.00 81.00 ;
        RECT 24.00 79.00 26.00 81.00 ;
        RECT 29.00 79.00 31.00 81.00 ;
        RECT 34.00 79.00 36.00 81.00 ;
        RECT 39.00 79.00 43.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 21.00 86.00 ;
        RECT 24.00 84.00 26.00 86.00 ;
        RECT 29.00 84.00 31.00 86.00 ;
        RECT 34.00 84.00 36.00 86.00 ;
        RECT 39.00 84.00 43.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 21.00 91.00 ;
        RECT 24.00 89.00 26.00 91.00 ;
        RECT 29.00 89.00 31.00 91.00 ;
        RECT 34.00 89.00 36.00 91.00 ;
        RECT 39.00 89.00 43.50 91.00 ;
        RECT 1.50 109.00 6.00 111.00 ;
        RECT 9.00 109.00 11.00 111.00 ;
        RECT 14.00 109.00 16.00 111.00 ;
        RECT 19.00 109.00 21.00 111.00 ;
        RECT 24.00 109.00 26.00 111.00 ;
        RECT 29.00 109.00 31.00 111.00 ;
        RECT 34.00 109.00 36.00 111.00 ;
        RECT 39.00 109.00 43.50 111.00 ;
        RECT 1.50 114.00 6.00 116.00 ;
        RECT 9.00 114.00 11.00 116.00 ;
        RECT 14.00 114.00 16.00 116.00 ;
        RECT 19.00 114.00 21.00 116.00 ;
        RECT 24.00 114.00 26.00 116.00 ;
        RECT 29.00 114.00 31.00 116.00 ;
        RECT 34.00 114.00 36.00 116.00 ;
        RECT 39.00 114.00 43.50 116.00 ;
        RECT 1.50 119.00 6.00 121.00 ;
        RECT 9.00 119.00 11.00 121.00 ;
        RECT 14.00 119.00 16.00 121.00 ;
        RECT 19.00 119.00 21.00 121.00 ;
        RECT 24.00 119.00 26.00 121.00 ;
        RECT 29.00 119.00 31.00 121.00 ;
        RECT 34.00 119.00 36.00 121.00 ;
        RECT 39.00 119.00 43.50 121.00 ;
        RECT 1.50 124.00 6.00 126.00 ;
        RECT 9.00 124.00 11.00 126.00 ;
        RECT 14.00 124.00 16.00 126.00 ;
        RECT 19.00 124.00 21.00 126.00 ;
        RECT 24.00 124.00 26.00 126.00 ;
        RECT 29.00 124.00 31.00 126.00 ;
        RECT 34.00 124.00 36.00 126.00 ;
        RECT 39.00 124.00 43.50 126.00 ;
        RECT 1.50 129.00 6.00 131.00 ;
        RECT 9.00 129.00 11.00 131.00 ;
        RECT 14.00 129.00 16.00 131.00 ;
        RECT 19.00 129.00 21.00 131.00 ;
        RECT 24.00 129.00 26.00 131.00 ;
        RECT 29.00 129.00 31.00 131.00 ;
        RECT 34.00 129.00 36.00 131.00 ;
        RECT 39.00 129.00 43.50 131.00 ;
        RECT 1.50 134.00 6.00 136.00 ;
        RECT 9.00 134.00 11.00 136.00 ;
        RECT 14.00 134.00 16.00 136.00 ;
        RECT 19.00 134.00 21.00 136.00 ;
        RECT 24.00 134.00 26.00 136.00 ;
        RECT 29.00 134.00 31.00 136.00 ;
        RECT 34.00 134.00 36.00 136.00 ;
        RECT 39.00 134.00 43.50 136.00 ;
        RECT 1.50 139.00 6.00 141.00 ;
        RECT 9.00 139.00 11.00 141.00 ;
        RECT 14.00 139.00 16.00 141.00 ;
        RECT 19.00 139.00 21.00 141.00 ;
        RECT 24.00 139.00 26.00 141.00 ;
        RECT 29.00 139.00 31.00 141.00 ;
        RECT 34.00 139.00 36.00 141.00 ;
        RECT 39.00 139.00 43.50 141.00 ;
        RECT 1.50 159.00 6.00 161.00 ;
        RECT 9.00 159.00 11.00 161.00 ;
        RECT 14.00 159.00 16.00 161.00 ;
        RECT 19.00 159.00 21.00 161.00 ;
        RECT 24.00 159.00 26.00 161.00 ;
        RECT 29.00 159.00 31.00 161.00 ;
        RECT 34.00 159.00 36.00 161.00 ;
        RECT 39.00 159.00 43.50 161.00 ;
        RECT 1.50 164.00 6.00 166.00 ;
        RECT 9.00 164.00 11.00 166.00 ;
        RECT 14.00 164.00 16.00 166.00 ;
        RECT 19.00 164.00 21.00 166.00 ;
        RECT 24.00 164.00 26.00 166.00 ;
        RECT 29.00 164.00 31.00 166.00 ;
        RECT 34.00 164.00 36.00 166.00 ;
        RECT 39.00 164.00 43.50 166.00 ;
        RECT 1.50 169.00 6.00 171.00 ;
        RECT 9.00 169.00 11.00 171.00 ;
        RECT 14.00 169.00 16.00 171.00 ;
        RECT 19.00 169.00 21.00 171.00 ;
        RECT 24.00 169.00 26.00 171.00 ;
        RECT 29.00 169.00 31.00 171.00 ;
        RECT 34.00 169.00 36.00 171.00 ;
        RECT 39.00 169.00 43.50 171.00 ;
        RECT 1.50 174.00 6.00 176.00 ;
        RECT 9.00 174.00 11.00 176.00 ;
        RECT 14.00 174.00 16.00 176.00 ;
        RECT 19.00 174.00 21.00 176.00 ;
        RECT 24.00 174.00 26.00 176.00 ;
        RECT 29.00 174.00 31.00 176.00 ;
        RECT 34.00 174.00 36.00 176.00 ;
        RECT 39.00 174.00 43.50 176.00 ;
        RECT 1.50 179.00 6.00 181.00 ;
        RECT 9.00 179.00 11.00 181.00 ;
        RECT 14.00 179.00 16.00 181.00 ;
        RECT 19.00 179.00 21.00 181.00 ;
        RECT 24.00 179.00 26.00 181.00 ;
        RECT 29.00 179.00 31.00 181.00 ;
        RECT 34.00 179.00 36.00 181.00 ;
        RECT 39.00 179.00 43.50 181.00 ;
        RECT 1.50 184.00 6.00 186.00 ;
        RECT 9.00 184.00 11.00 186.00 ;
        RECT 14.00 184.00 16.00 186.00 ;
        RECT 19.00 184.00 21.00 186.00 ;
        RECT 24.00 184.00 26.00 186.00 ;
        RECT 29.00 184.00 31.00 186.00 ;
        RECT 34.00 184.00 36.00 186.00 ;
        RECT 39.00 184.00 43.50 186.00 ;
        RECT 1.50 189.00 6.00 191.00 ;
        RECT 9.00 189.00 11.00 191.00 ;
        RECT 14.00 189.00 16.00 191.00 ;
        RECT 19.00 189.00 21.00 191.00 ;
        RECT 24.00 189.00 26.00 191.00 ;
        RECT 29.00 189.00 31.00 191.00 ;
        RECT 34.00 189.00 36.00 191.00 ;
        RECT 39.00 189.00 43.50 191.00 ;
        LAYER L_ALU2 ;
        RECT 26.00 39.00 40.00 41.00 ;
        RECT 8.00 14.00 26.00 16.00 ;
        RECT 26.00 159.00 40.00 161.00 ;
        RECT 8.00 184.00 26.00 186.00 ;
        RECT 26.00 39.00 40.00 41.00 ;
        RECT 8.00 14.00 26.00 16.00 ;
        RECT 8.00 184.00 26.00 186.00 ;
        RECT 26.00 159.00 40.00 161.00 ;
        RECT 4.00 99.00 16.00 101.00 ;
        RECT 4.00 -1.00 16.00 1.00 ;
        RECT 4.00 199.00 16.00 201.00 ;
    END
END rf_inmux_buf_4


MACRO rf_inmux_mem
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN dinx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END dinx
    PIN sel1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 29.00 26.00 31.00 ;
        END
    END sel1
    PIN sel0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 29.00 36.00 31.00 ;
        END
    END sel0
    PIN datain0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END datain0
    PIN datain1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END datain1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 10.00 6.00 10.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 43.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 43.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 43.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 43.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 43.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 43.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 43.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 24.00 29.00 36.00 31.00 ;
        RECT 4.00 -1.00 16.00 1.00 ;
    END
END rf_inmux_mem


MACRO rf_mid_buf_2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN write
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END write
    PIN read
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END read
    PIN nck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 89.00 26.00 91.00 ;
        END
    END nck
    PIN selr
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 79.00 11.00 81.00 ;
        END
    END selr
    PIN selw
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 84.00 16.00 86.00 ;
        END
    END selw
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 22.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 22.00 97.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 23.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 23.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 23.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 23.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 23.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 23.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 23.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 23.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 23.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 23.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 23.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 23.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 23.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 23.50 91.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 14.00 21.00 16.00 ;
        RECT 4.00 39.00 21.00 41.00 ;
        RECT 4.00 59.00 21.00 61.00 ;
    END
END rf_mid_buf_2


MACRO rf_mid_buf_4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 200.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN read
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 184.00 6.00 186.00 ;
            RECT 4.00 179.00 6.00 181.00 ;
            RECT 4.00 174.00 6.00 176.00 ;
            RECT 4.00 169.00 6.00 171.00 ;
            RECT 4.00 164.00 6.00 166.00 ;
            RECT 4.00 159.00 6.00 161.00 ;
            RECT 4.00 154.00 6.00 156.00 ;
            RECT 4.00 149.00 6.00 151.00 ;
            RECT 4.00 144.00 6.00 146.00 ;
            RECT 4.00 139.00 6.00 141.00 ;
        END
    END read
    PIN write
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END write
    PIN nck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 9.00 89.00 11.00 91.00 ;
            RECT 4.00 89.00 6.00 91.00 ;
            RECT -1.00 89.00 1.00 91.00 ;
        END
    END nck
    PIN selw
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 84.00 16.00 86.00 ;
        END
    END selw
    PIN selr
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 114.00 11.00 116.00 ;
        END
    END selr
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 22.00 53.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 147.00 22.00 147.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 153.00 22.00 153.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 22.00 97.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 103.00 22.00 103.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 197.00 22.00 197.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 23.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 23.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 23.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 23.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 23.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 23.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 23.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 23.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 23.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 23.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 23.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 23.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 23.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 23.50 91.00 ;
        RECT 1.50 109.00 6.00 111.00 ;
        RECT 9.00 109.00 11.00 111.00 ;
        RECT 14.00 109.00 16.00 111.00 ;
        RECT 19.00 109.00 23.50 111.00 ;
        RECT 1.50 114.00 6.00 116.00 ;
        RECT 9.00 114.00 11.00 116.00 ;
        RECT 14.00 114.00 16.00 116.00 ;
        RECT 19.00 114.00 23.50 116.00 ;
        RECT 1.50 119.00 6.00 121.00 ;
        RECT 9.00 119.00 11.00 121.00 ;
        RECT 14.00 119.00 16.00 121.00 ;
        RECT 19.00 119.00 23.50 121.00 ;
        RECT 1.50 124.00 6.00 126.00 ;
        RECT 9.00 124.00 11.00 126.00 ;
        RECT 14.00 124.00 16.00 126.00 ;
        RECT 19.00 124.00 23.50 126.00 ;
        RECT 1.50 129.00 6.00 131.00 ;
        RECT 9.00 129.00 11.00 131.00 ;
        RECT 14.00 129.00 16.00 131.00 ;
        RECT 19.00 129.00 23.50 131.00 ;
        RECT 1.50 134.00 6.00 136.00 ;
        RECT 9.00 134.00 11.00 136.00 ;
        RECT 14.00 134.00 16.00 136.00 ;
        RECT 19.00 134.00 23.50 136.00 ;
        RECT 1.50 139.00 6.00 141.00 ;
        RECT 9.00 139.00 11.00 141.00 ;
        RECT 14.00 139.00 16.00 141.00 ;
        RECT 19.00 139.00 23.50 141.00 ;
        RECT 1.50 159.00 6.00 161.00 ;
        RECT 9.00 159.00 11.00 161.00 ;
        RECT 14.00 159.00 16.00 161.00 ;
        RECT 19.00 159.00 23.50 161.00 ;
        RECT 1.50 164.00 6.00 166.00 ;
        RECT 9.00 164.00 11.00 166.00 ;
        RECT 14.00 164.00 16.00 166.00 ;
        RECT 19.00 164.00 23.50 166.00 ;
        RECT 1.50 169.00 6.00 171.00 ;
        RECT 9.00 169.00 11.00 171.00 ;
        RECT 14.00 169.00 16.00 171.00 ;
        RECT 19.00 169.00 23.50 171.00 ;
        RECT 1.50 174.00 6.00 176.00 ;
        RECT 9.00 174.00 11.00 176.00 ;
        RECT 14.00 174.00 16.00 176.00 ;
        RECT 19.00 174.00 23.50 176.00 ;
        RECT 1.50 179.00 6.00 181.00 ;
        RECT 9.00 179.00 11.00 181.00 ;
        RECT 14.00 179.00 16.00 181.00 ;
        RECT 19.00 179.00 23.50 181.00 ;
        RECT 1.50 184.00 6.00 186.00 ;
        RECT 9.00 184.00 11.00 186.00 ;
        RECT 14.00 184.00 16.00 186.00 ;
        RECT 19.00 184.00 23.50 186.00 ;
        RECT 1.50 189.00 6.00 191.00 ;
        RECT 9.00 189.00 11.00 191.00 ;
        RECT 14.00 189.00 16.00 191.00 ;
        RECT 19.00 189.00 23.50 191.00 ;
        LAYER L_ALU2 ;
        RECT -1.00 14.00 26.00 16.00 ;
        RECT -1.00 39.00 26.00 41.00 ;
        RECT -1.00 59.00 26.00 61.00 ;
        RECT -1.00 139.00 26.00 141.00 ;
        RECT -1.00 159.00 26.00 161.00 ;
        RECT -1.00 184.00 26.00 186.00 ;
    END
END rf_mid_buf_4


MACRO rf_mid_mem
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN rbus
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 24.00 26.00 26.00 ;
        END
    END rbus
    PIN read
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END read
    PIN write
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END write
    PIN dinx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END dinx
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 23.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 23.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 23.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 23.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 23.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 23.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 23.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 29.00 16.00 31.00 ;
        RECT 4.00 29.00 16.00 31.00 ;
        RECT 19.00 14.00 26.00 16.00 ;
    END
END rf_mid_mem


MACRO rf_mid_mem_r0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN rbus
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 24.00 26.00 26.00 ;
        END
    END rbus
    PIN dinx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END dinx
    PIN write
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END write
    PIN read
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END read
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 23.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 23.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 23.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 23.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 23.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 23.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 23.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 29.00 16.00 31.00 ;
        RECT 4.00 29.00 16.00 31.00 ;
        RECT 19.00 14.00 26.00 16.00 ;
    END
END rf_mid_mem_r0


MACRO rf_out_buf_2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      55.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN xcks
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 59.00 16.00 61.00 ;
            RECT 14.00 54.00 16.00 56.00 ;
            RECT 14.00 49.00 16.00 51.00 ;
            RECT 14.00 44.00 16.00 46.00 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END xcks
    PIN nck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 89.00 16.00 91.00 ;
        END
    END nck
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 52.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 52.00 53.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 45.00 6.00 45.00 94.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 52.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 52.00 97.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 53.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 53.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 53.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 53.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 53.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 53.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 53.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 21.00 61.00 ;
        RECT 24.00 59.00 26.00 61.00 ;
        RECT 29.00 59.00 31.00 61.00 ;
        RECT 34.00 59.00 36.00 61.00 ;
        RECT 39.00 59.00 41.00 61.00 ;
        RECT 44.00 59.00 46.00 61.00 ;
        RECT 49.00 59.00 53.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 26.00 66.00 ;
        RECT 29.00 64.00 31.00 66.00 ;
        RECT 34.00 64.00 36.00 66.00 ;
        RECT 39.00 64.00 41.00 66.00 ;
        RECT 44.00 64.00 46.00 66.00 ;
        RECT 49.00 64.00 53.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 21.00 71.00 ;
        RECT 24.00 69.00 26.00 71.00 ;
        RECT 29.00 69.00 31.00 71.00 ;
        RECT 34.00 69.00 36.00 71.00 ;
        RECT 39.00 69.00 41.00 71.00 ;
        RECT 44.00 69.00 46.00 71.00 ;
        RECT 49.00 69.00 53.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 21.00 76.00 ;
        RECT 24.00 74.00 26.00 76.00 ;
        RECT 29.00 74.00 31.00 76.00 ;
        RECT 34.00 74.00 36.00 76.00 ;
        RECT 39.00 74.00 41.00 76.00 ;
        RECT 44.00 74.00 46.00 76.00 ;
        RECT 49.00 74.00 53.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 21.00 81.00 ;
        RECT 24.00 79.00 26.00 81.00 ;
        RECT 29.00 79.00 31.00 81.00 ;
        RECT 34.00 79.00 36.00 81.00 ;
        RECT 39.00 79.00 41.00 81.00 ;
        RECT 44.00 79.00 46.00 81.00 ;
        RECT 49.00 79.00 53.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 21.00 86.00 ;
        RECT 24.00 84.00 26.00 86.00 ;
        RECT 29.00 84.00 31.00 86.00 ;
        RECT 34.00 84.00 36.00 86.00 ;
        RECT 39.00 84.00 41.00 86.00 ;
        RECT 44.00 84.00 46.00 86.00 ;
        RECT 49.00 84.00 53.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 21.00 91.00 ;
        RECT 24.00 89.00 26.00 91.00 ;
        RECT 29.00 89.00 31.00 91.00 ;
        RECT 34.00 89.00 36.00 91.00 ;
        RECT 39.00 89.00 41.00 91.00 ;
        RECT 44.00 89.00 46.00 91.00 ;
        RECT 49.00 89.00 53.50 91.00 ;
        LAYER L_ALU2 ;
        RECT 39.00 49.00 51.00 51.00 ;
        RECT 9.00 14.00 21.00 16.00 ;
        RECT 9.00 39.00 21.00 41.00 ;
        RECT 9.00 59.00 21.00 61.00 ;
    END
END rf_out_buf_2


MACRO rf_out_buf_4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      55.00 BY 200.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN xcks
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 184.00 16.00 186.00 ;
            RECT 14.00 179.00 16.00 181.00 ;
            RECT 14.00 174.00 16.00 176.00 ;
            RECT 14.00 169.00 16.00 171.00 ;
            RECT 14.00 164.00 16.00 166.00 ;
            RECT 14.00 159.00 16.00 161.00 ;
            RECT 14.00 154.00 16.00 156.00 ;
            RECT 14.00 149.00 16.00 151.00 ;
            RECT 14.00 144.00 16.00 146.00 ;
            RECT 14.00 139.00 16.00 141.00 ;
            RECT 14.00 134.00 16.00 136.00 ;
            RECT 14.00 129.00 16.00 131.00 ;
            RECT 14.00 124.00 16.00 126.00 ;
            RECT 14.00 119.00 16.00 121.00 ;
            RECT 14.00 114.00 16.00 116.00 ;
            RECT 14.00 109.00 16.00 111.00 ;
            RECT 14.00 104.00 16.00 106.00 ;
            RECT 14.00 99.00 16.00 101.00 ;
            RECT 14.00 94.00 16.00 96.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 14.00 79.00 16.00 81.00 ;
            RECT 14.00 74.00 16.00 76.00 ;
            RECT 14.00 69.00 16.00 71.00 ;
            RECT 14.00 64.00 16.00 66.00 ;
            RECT 14.00 59.00 16.00 61.00 ;
            RECT 14.00 54.00 16.00 56.00 ;
            RECT 14.00 49.00 16.00 51.00 ;
            RECT 14.00 44.00 16.00 46.00 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END xcks
    PIN nck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 89.00 16.00 91.00 ;
        END
    END nck
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 52.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 52.00 53.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 147.00 52.00 147.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 153.00 52.00 153.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 45.00 6.00 45.00 194.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 52.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 52.00 97.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 103.00 52.00 103.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 197.00 52.00 197.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 53.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 53.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 53.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 53.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 53.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 53.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 53.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 21.00 61.00 ;
        RECT 24.00 59.00 26.00 61.00 ;
        RECT 29.00 59.00 31.00 61.00 ;
        RECT 34.00 59.00 36.00 61.00 ;
        RECT 39.00 59.00 41.00 61.00 ;
        RECT 44.00 59.00 46.00 61.00 ;
        RECT 49.00 59.00 53.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 26.00 66.00 ;
        RECT 29.00 64.00 31.00 66.00 ;
        RECT 34.00 64.00 36.00 66.00 ;
        RECT 39.00 64.00 41.00 66.00 ;
        RECT 44.00 64.00 46.00 66.00 ;
        RECT 49.00 64.00 53.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 21.00 71.00 ;
        RECT 24.00 69.00 26.00 71.00 ;
        RECT 29.00 69.00 31.00 71.00 ;
        RECT 34.00 69.00 36.00 71.00 ;
        RECT 39.00 69.00 41.00 71.00 ;
        RECT 44.00 69.00 46.00 71.00 ;
        RECT 49.00 69.00 53.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 21.00 76.00 ;
        RECT 24.00 74.00 26.00 76.00 ;
        RECT 29.00 74.00 31.00 76.00 ;
        RECT 34.00 74.00 36.00 76.00 ;
        RECT 39.00 74.00 41.00 76.00 ;
        RECT 44.00 74.00 46.00 76.00 ;
        RECT 49.00 74.00 53.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 21.00 81.00 ;
        RECT 24.00 79.00 26.00 81.00 ;
        RECT 29.00 79.00 31.00 81.00 ;
        RECT 34.00 79.00 36.00 81.00 ;
        RECT 39.00 79.00 41.00 81.00 ;
        RECT 44.00 79.00 46.00 81.00 ;
        RECT 49.00 79.00 53.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 21.00 86.00 ;
        RECT 24.00 84.00 26.00 86.00 ;
        RECT 29.00 84.00 31.00 86.00 ;
        RECT 34.00 84.00 36.00 86.00 ;
        RECT 39.00 84.00 41.00 86.00 ;
        RECT 44.00 84.00 46.00 86.00 ;
        RECT 49.00 84.00 53.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 21.00 91.00 ;
        RECT 24.00 89.00 26.00 91.00 ;
        RECT 29.00 89.00 31.00 91.00 ;
        RECT 34.00 89.00 36.00 91.00 ;
        RECT 39.00 89.00 41.00 91.00 ;
        RECT 44.00 89.00 46.00 91.00 ;
        RECT 49.00 89.00 53.50 91.00 ;
        RECT 1.50 109.00 6.00 111.00 ;
        RECT 9.00 109.00 11.00 111.00 ;
        RECT 14.00 109.00 16.00 111.00 ;
        RECT 19.00 109.00 21.00 111.00 ;
        RECT 24.00 109.00 26.00 111.00 ;
        RECT 29.00 109.00 31.00 111.00 ;
        RECT 34.00 109.00 36.00 111.00 ;
        RECT 39.00 109.00 41.00 111.00 ;
        RECT 44.00 109.00 46.00 111.00 ;
        RECT 49.00 109.00 53.50 111.00 ;
        RECT 1.50 114.00 6.00 116.00 ;
        RECT 9.00 114.00 11.00 116.00 ;
        RECT 14.00 114.00 16.00 116.00 ;
        RECT 19.00 114.00 21.00 116.00 ;
        RECT 24.00 114.00 26.00 116.00 ;
        RECT 29.00 114.00 31.00 116.00 ;
        RECT 34.00 114.00 36.00 116.00 ;
        RECT 39.00 114.00 41.00 116.00 ;
        RECT 44.00 114.00 46.00 116.00 ;
        RECT 49.00 114.00 53.50 116.00 ;
        RECT 1.50 119.00 6.00 121.00 ;
        RECT 9.00 119.00 11.00 121.00 ;
        RECT 14.00 119.00 16.00 121.00 ;
        RECT 19.00 119.00 21.00 121.00 ;
        RECT 24.00 119.00 26.00 121.00 ;
        RECT 29.00 119.00 31.00 121.00 ;
        RECT 34.00 119.00 36.00 121.00 ;
        RECT 39.00 119.00 41.00 121.00 ;
        RECT 44.00 119.00 46.00 121.00 ;
        RECT 49.00 119.00 53.50 121.00 ;
        RECT 1.50 124.00 6.00 126.00 ;
        RECT 9.00 124.00 11.00 126.00 ;
        RECT 14.00 124.00 16.00 126.00 ;
        RECT 19.00 124.00 21.00 126.00 ;
        RECT 24.00 124.00 26.00 126.00 ;
        RECT 29.00 124.00 31.00 126.00 ;
        RECT 34.00 124.00 36.00 126.00 ;
        RECT 39.00 124.00 41.00 126.00 ;
        RECT 44.00 124.00 46.00 126.00 ;
        RECT 49.00 124.00 53.50 126.00 ;
        RECT 1.50 129.00 6.00 131.00 ;
        RECT 9.00 129.00 11.00 131.00 ;
        RECT 14.00 129.00 16.00 131.00 ;
        RECT 19.00 129.00 21.00 131.00 ;
        RECT 24.00 129.00 26.00 131.00 ;
        RECT 29.00 129.00 31.00 131.00 ;
        RECT 34.00 129.00 36.00 131.00 ;
        RECT 39.00 129.00 41.00 131.00 ;
        RECT 44.00 129.00 46.00 131.00 ;
        RECT 49.00 129.00 53.50 131.00 ;
        RECT 1.50 134.00 6.00 136.00 ;
        RECT 9.00 134.00 11.00 136.00 ;
        RECT 14.00 134.00 16.00 136.00 ;
        RECT 19.00 134.00 21.00 136.00 ;
        RECT 24.00 134.00 26.00 136.00 ;
        RECT 29.00 134.00 31.00 136.00 ;
        RECT 34.00 134.00 36.00 136.00 ;
        RECT 39.00 134.00 41.00 136.00 ;
        RECT 44.00 134.00 46.00 136.00 ;
        RECT 49.00 134.00 53.50 136.00 ;
        RECT 1.50 139.00 6.00 141.00 ;
        RECT 9.00 139.00 11.00 141.00 ;
        RECT 14.00 139.00 16.00 141.00 ;
        RECT 19.00 139.00 21.00 141.00 ;
        RECT 24.00 139.00 26.00 141.00 ;
        RECT 29.00 139.00 31.00 141.00 ;
        RECT 34.00 139.00 36.00 141.00 ;
        RECT 39.00 139.00 41.00 141.00 ;
        RECT 44.00 139.00 46.00 141.00 ;
        RECT 49.00 139.00 53.50 141.00 ;
        RECT 1.50 159.00 6.00 161.00 ;
        RECT 9.00 159.00 11.00 161.00 ;
        RECT 14.00 159.00 16.00 161.00 ;
        RECT 19.00 159.00 21.00 161.00 ;
        RECT 24.00 159.00 26.00 161.00 ;
        RECT 29.00 159.00 31.00 161.00 ;
        RECT 34.00 159.00 36.00 161.00 ;
        RECT 39.00 159.00 41.00 161.00 ;
        RECT 44.00 159.00 46.00 161.00 ;
        RECT 49.00 159.00 53.50 161.00 ;
        RECT 1.50 164.00 6.00 166.00 ;
        RECT 9.00 164.00 11.00 166.00 ;
        RECT 14.00 164.00 16.00 166.00 ;
        RECT 19.00 164.00 21.00 166.00 ;
        RECT 24.00 164.00 26.00 166.00 ;
        RECT 29.00 164.00 31.00 166.00 ;
        RECT 34.00 164.00 36.00 166.00 ;
        RECT 39.00 164.00 41.00 166.00 ;
        RECT 44.00 164.00 46.00 166.00 ;
        RECT 49.00 164.00 53.50 166.00 ;
        RECT 1.50 169.00 6.00 171.00 ;
        RECT 9.00 169.00 11.00 171.00 ;
        RECT 14.00 169.00 16.00 171.00 ;
        RECT 19.00 169.00 21.00 171.00 ;
        RECT 24.00 169.00 26.00 171.00 ;
        RECT 29.00 169.00 31.00 171.00 ;
        RECT 34.00 169.00 36.00 171.00 ;
        RECT 39.00 169.00 41.00 171.00 ;
        RECT 44.00 169.00 46.00 171.00 ;
        RECT 49.00 169.00 53.50 171.00 ;
        RECT 1.50 174.00 6.00 176.00 ;
        RECT 9.00 174.00 11.00 176.00 ;
        RECT 14.00 174.00 16.00 176.00 ;
        RECT 19.00 174.00 21.00 176.00 ;
        RECT 24.00 174.00 26.00 176.00 ;
        RECT 29.00 174.00 31.00 176.00 ;
        RECT 34.00 174.00 36.00 176.00 ;
        RECT 39.00 174.00 41.00 176.00 ;
        RECT 44.00 174.00 46.00 176.00 ;
        RECT 49.00 174.00 53.50 176.00 ;
        RECT 1.50 179.00 6.00 181.00 ;
        RECT 9.00 179.00 11.00 181.00 ;
        RECT 14.00 179.00 16.00 181.00 ;
        RECT 19.00 179.00 21.00 181.00 ;
        RECT 24.00 179.00 26.00 181.00 ;
        RECT 29.00 179.00 31.00 181.00 ;
        RECT 34.00 179.00 36.00 181.00 ;
        RECT 39.00 179.00 41.00 181.00 ;
        RECT 44.00 179.00 46.00 181.00 ;
        RECT 49.00 179.00 53.50 181.00 ;
        RECT 1.50 184.00 6.00 186.00 ;
        RECT 9.00 184.00 11.00 186.00 ;
        RECT 14.00 184.00 16.00 186.00 ;
        RECT 19.00 184.00 21.00 186.00 ;
        RECT 24.00 184.00 26.00 186.00 ;
        RECT 29.00 184.00 31.00 186.00 ;
        RECT 34.00 184.00 36.00 186.00 ;
        RECT 39.00 184.00 41.00 186.00 ;
        RECT 44.00 184.00 46.00 186.00 ;
        RECT 49.00 184.00 53.50 186.00 ;
        RECT 1.50 189.00 6.00 191.00 ;
        RECT 9.00 189.00 11.00 191.00 ;
        RECT 14.00 189.00 16.00 191.00 ;
        RECT 19.00 189.00 21.00 191.00 ;
        RECT 24.00 189.00 26.00 191.00 ;
        RECT 29.00 189.00 31.00 191.00 ;
        RECT 34.00 189.00 36.00 191.00 ;
        RECT 39.00 189.00 41.00 191.00 ;
        RECT 44.00 189.00 46.00 191.00 ;
        RECT 49.00 189.00 53.50 191.00 ;
        LAYER L_ALU2 ;
        RECT 39.00 149.00 51.00 151.00 ;
        RECT 39.00 49.00 51.00 51.00 ;
        RECT 9.00 14.00 21.00 16.00 ;
        RECT 9.00 39.00 21.00 41.00 ;
        RECT 9.00 59.00 21.00 61.00 ;
        RECT 9.00 139.00 21.00 141.00 ;
        RECT 9.00 159.00 21.00 161.00 ;
        RECT 9.00 184.00 21.00 186.00 ;
    END
END rf_out_buf_4


MACRO rf_out_mem
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      55.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN dataout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 39.00 46.00 41.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
        END
    END dataout
    PIN rbus
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 4.00 24.00 6.00 26.00 ;
        END
    END rbus
    PIN xcks
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END xcks
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 52.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 45.00 6.00 45.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 52.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 53.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 53.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 53.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 53.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 53.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 53.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 53.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 39.00 49.00 51.00 51.00 ;
        RECT 14.00 24.00 24.00 26.00 ;
        RECT 14.00 24.00 26.00 26.00 ;
    END
END rf_out_mem


END LIBRARY
