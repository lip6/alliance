
VERSION             5.2 ;
NAMESCASESENSITIVE  ON ;
BUSBITCHARS         "()" ;
DIVIDERCHAR         "." ;


MACRO a2_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
    END
END a2_x2


MACRO a2_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END a2_x4


MACRO a3_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END a3_x2


MACRO a3_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END a3_x4


MACRO a4_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END q
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i3
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i2
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END a4_x2


MACRO a4_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END q
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i3
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i2
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END a4_x4


MACRO an12_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
    END
END an12_x1


MACRO an12_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END an12_x4


MACRO ao22_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END q
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END ao22_x2


MACRO ao22_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END ao22_x4


MACRO ao2o22_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 43.50 41.00 ;
    END
END ao2o22_x2


MACRO ao2o22_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END ao2o22_x4


MACRO buf_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      20.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 17.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 17.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 18.50 41.00 ;
    END
END buf_x2


MACRO buf_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
    END
END buf_x4


MACRO buf_x8
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END buf_x8


MACRO fulladder_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      100.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN cout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            LAYER L_ALU1 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END cout
    PIN sout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END sout
    PIN cin1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END cin1
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END a2
    PIN b2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END b2
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
        END
    END a3
    PIN b3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 64.00 29.00 66.00 31.00 ;
            RECT 64.00 24.00 66.00 26.00 ;
            RECT 64.00 19.00 66.00 21.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
        END
    END b3
    PIN cin2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
        END
    END cin2
    PIN cin3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 84.00 29.00 86.00 31.00 ;
            RECT 84.00 24.00 86.00 26.00 ;
            RECT 84.00 19.00 86.00 21.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
        END
    END cin3
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a1
    PIN b1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END b1
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 89.00 34.00 91.00 36.00 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
        END
    END a4
    PIN b4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
        END
    END b4
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 97.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 97.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 98.50 41.00 ;
    END
END fulladder_x2


MACRO fulladder_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      105.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN sout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
        END
    END sout
    PIN cout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
        END
    END cout
    PIN a1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END a1
    PIN b1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END b1
    PIN cin1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END cin1
    PIN a2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END a2
    PIN b2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END b2
    PIN b4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
            RECT 99.00 14.00 101.00 16.00 ;
        END
    END b4
    PIN a4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 94.00 34.00 96.00 36.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 94.00 19.00 96.00 21.00 ;
            RECT 94.00 14.00 96.00 16.00 ;
        END
    END a4
    PIN cin3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 89.00 29.00 91.00 31.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 89.00 19.00 91.00 21.00 ;
            RECT 89.00 14.00 91.00 16.00 ;
        END
    END cin3
    PIN b3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
        END
    END b3
    PIN cin2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 74.00 29.00 76.00 31.00 ;
            RECT 74.00 24.00 76.00 26.00 ;
            RECT 74.00 19.00 76.00 21.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
        END
    END cin2
    PIN a3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 64.00 29.00 66.00 31.00 ;
            RECT 64.00 24.00 66.00 26.00 ;
            RECT 64.00 19.00 66.00 21.00 ;
        END
    END a3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 102.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 102.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 103.50 41.00 ;
    END
END fulladder_x4


MACRO halfadder_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      80.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN sout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 74.00 39.00 76.00 41.00 ;
            RECT 74.00 34.00 76.00 36.00 ;
            RECT 74.00 29.00 76.00 31.00 ;
            RECT 74.00 24.00 76.00 26.00 ;
            RECT 74.00 19.00 76.00 21.00 ;
            RECT 74.00 14.00 76.00 16.00 ;
            RECT 74.00 9.00 76.00 11.00 ;
        END
    END sout
    PIN cout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END cout
    PIN b
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
        END
    END b
    PIN a
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END a
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 77.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 77.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 78.50 41.00 ;
    END
END halfadder_x2


MACRO halfadder_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      90.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN sout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END sout
    PIN cout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END cout
    PIN b
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END b
    PIN a
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END a
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 87.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 87.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 88.50 41.00 ;
    END
END halfadder_x4


MACRO inv_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      15.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 12.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 12.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 13.50 41.00 ;
    END
END inv_x1


MACRO inv_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      15.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 12.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 12.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 13.50 41.00 ;
    END
END inv_x2


MACRO inv_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      20.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 17.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 17.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 18.50 41.00 ;
    END
END inv_x4


MACRO inv_x8
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END inv_x8


MACRO mx2_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END q
    PIN cmd
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END cmd
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 43.50 41.00 ;
    END
END mx2_x2


MACRO mx2_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END q
    PIN cmd
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END cmd
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END mx2_x4


MACRO mx3_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      65.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            LAYER L_ALU1 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
        END
    END q
    PIN cmd1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END cmd1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 24.00 26.00 26.00 ;
        END
    END i1
    PIN cmd0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END cmd0
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 19.00 41.00 21.00 ;
            LAYER L_ALU1 ;
            RECT 44.00 24.00 46.00 26.00 ;
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 62.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 62.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 63.50 41.00 ;
    END
END mx3_x2


MACRO mx3_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      70.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 64.00 19.00 66.00 21.00 ;
            LAYER L_ALU1 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
            LAYER L_ALU1 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
        END
    END q
    PIN cmd0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END cmd0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 24.00 26.00 26.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END i2
    PIN cmd1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END cmd1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 19.00 41.00 21.00 ;
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            LAYER L_ALU1 ;
            RECT 44.00 24.00 46.00 26.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 67.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 67.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 68.50 41.00 ;
    END
END mx3_x4


MACRO na2_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      20.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 17.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 17.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 18.50 41.00 ;
    END
END na2_x1


MACRO na2_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END na2_x4


MACRO na3_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
    END
END na3_x1


MACRO na3_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END nq
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END na3_x4


MACRO na4_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END na4_x1


MACRO na4_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nq
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END i3
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END na4_x4


MACRO nao22_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END nao22_x1


MACRO nao22_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END nq
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 14.00 26.00 16.00 ;
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END nao22_x4


MACRO nao2o22_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i1
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END nao2o22_x1


MACRO nao2o22_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      55.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 39.00 46.00 41.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i1
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 52.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 52.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 53.50 41.00 ;
    END
END nao2o22_x4


MACRO nmx2_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            LAYER L_ALU1 ;
            RECT 19.00 9.00 21.00 11.00 ;
            LAYER L_ALU1 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i0
    PIN cmd
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END cmd
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END nmx2_x1


MACRO nmx2_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      60.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i0
    PIN cmd
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END cmd
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 57.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 57.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 58.50 41.00 ;
    END
END nmx2_x4


MACRO nmx3_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      60.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            LAYER L_ALU1 ;
            RECT 44.00 24.00 46.00 26.00 ;
            LAYER L_ALU1 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END i0
    PIN cmd1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END cmd1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 24.00 26.00 26.00 ;
        END
    END i1
    PIN cmd0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END cmd0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 57.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 57.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 58.50 41.00 ;
    END
END nmx3_x1


MACRO nmx3_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      75.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
        END
    END nq
    PIN cmd0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END cmd0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 24.00 26.00 26.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END i2
    PIN cmd1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END cmd1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 19.00 41.00 21.00 ;
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            LAYER L_ALU1 ;
            RECT 44.00 24.00 46.00 26.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 72.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 72.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 73.50 41.00 ;
    END
END nmx3_x4


MACRO no2_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      20.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 17.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 17.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 18.50 41.00 ;
    END
END no2_x1


MACRO no2_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END no2_x4


MACRO no3_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END nq
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
    END
END no3_x1


MACRO no3_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END nq
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END no3_x4


MACRO no4_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END nq
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i3
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END no4_x1


MACRO no4_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 39.00 36.00 41.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END nq
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i3
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END no4_x4


MACRO noa22_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END noa22_x1


MACRO noa22_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END noa22_x4


MACRO noa2a22_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nq
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i3
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END noa2a22_x1


MACRO noa2a22_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      55.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 39.00 46.00 41.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 52.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 52.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 53.50 41.00 ;
    END
END noa2a22_x4


MACRO noa2a2a23_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END nq
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i5
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i3
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i1
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i4
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END noa2a2a23_x1


MACRO noa2a2a23_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      65.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i0
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i4
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i3
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i5
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 62.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 62.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 63.50 41.00 ;
    END
END noa2a2a23_x4


MACRO noa2a2a2a24_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      70.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END i3
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i4
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i5
    PIN i6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i6
    PIN i7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i7
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 67.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 67.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 68.50 41.00 ;
    END
END noa2a2a2a24_x1


MACRO noa2a2a2a24_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      85.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
        END
    END nq
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END i3
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i4
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i5
    PIN i6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i6
    PIN i7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i7
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 64.00 34.00 66.00 36.00 ;
            RECT 64.00 29.00 66.00 31.00 ;
            RECT 64.00 24.00 66.00 26.00 ;
            RECT 64.00 19.00 66.00 21.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 82.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 82.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 83.50 41.00 ;
    END
END noa2a2a2a24_x4


MACRO noa2ao222_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            LAYER L_ALU1 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nq
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i4
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END noa2ao222_x1


MACRO noa2ao222_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      60.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i4
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 57.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 57.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 58.50 41.00 ;
    END
END noa2ao222_x4


MACRO noa3ao322_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i2
    PIN i6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i6
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i3
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END i4
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i5
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 43.50 41.00 ;
    END
END noa3ao322_x1


MACRO noa3ao322_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      65.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i0
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
        END
    END i3
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
        END
    END i5
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
        END
    END i4
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END i2
    PIN i6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END i6
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 62.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 62.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 63.50 41.00 ;
    END
END noa3ao322_x4


MACRO nts_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nq
    PIN cmd
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END cmd
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END nts_x1


MACRO nts_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i
    PIN cmd
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END cmd
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END nts_x2


MACRO nxr2_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 39.00 36.00 41.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 43.50 41.00 ;
    END
END nxr2_x1


MACRO nxr2_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      60.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 39.00 36.00 41.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 57.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 57.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 58.50 41.00 ;
    END
END nxr2_x4


MACRO o2_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
    END
END o2_x2


MACRO o2_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END o2_x4


MACRO o3_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END q
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END o3_x2


MACRO o3_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END o3_x4


MACRO o4_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END o4_x2


MACRO o4_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
        END
    END q
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i3
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END o4_x4


MACRO oa22_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
    END
END oa22_x2


MACRO oa22_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END q
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END oa22_x4


MACRO oa2a22_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END q
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 43.50 41.00 ;
    END
END oa2a22_x2


MACRO oa2a22_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
            RECT 39.00 9.00 41.00 11.00 ;
        END
    END q
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END oa2a22_x4


MACRO oa2a2a23_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      60.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 39.00 56.00 41.00 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i1
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i4
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i5
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 57.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 57.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 58.50 41.00 ;
    END
END oa2a2a23_x2


MACRO oa2a2a23_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      65.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 39.00 56.00 41.00 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
            RECT 54.00 9.00 56.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
        END
    END i0
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i4
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i3
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i5
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 62.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 62.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 63.50 41.00 ;
    END
END oa2a2a23_x4


MACRO oa2a2a2a24_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      75.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END q
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END i3
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i4
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i5
    PIN i6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i6
    PIN i7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i7
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 64.00 34.00 66.00 36.00 ;
            RECT 64.00 29.00 66.00 31.00 ;
            RECT 64.00 24.00 66.00 26.00 ;
            RECT 64.00 19.00 66.00 21.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 72.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 72.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 73.50 41.00 ;
    END
END oa2a2a2a24_x2


MACRO oa2a2a2a24_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      80.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 69.00 39.00 71.00 41.00 ;
            RECT 69.00 34.00 71.00 36.00 ;
            RECT 69.00 29.00 71.00 31.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 69.00 19.00 71.00 21.00 ;
            RECT 69.00 14.00 71.00 16.00 ;
            RECT 69.00 9.00 71.00 11.00 ;
        END
    END q
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END i3
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i4
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i5
    PIN i6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i6
    PIN i7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i7
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 64.00 34.00 66.00 36.00 ;
            RECT 64.00 29.00 66.00 31.00 ;
            RECT 64.00 24.00 66.00 26.00 ;
            RECT 64.00 19.00 66.00 21.00 ;
            RECT 64.00 14.00 66.00 16.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 77.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 77.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 78.50 41.00 ;
    END
END oa2a2a2a24_x4


MACRO oa2ao222_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 39.00 46.00 41.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i4
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END oa2ao222_x2


MACRO oa2ao222_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      55.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 39.00 46.00 41.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
        END
    END q
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i2
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i4
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 52.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 52.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 53.50 41.00 ;
    END
END oa2ao222_x4


MACRO oa3ao322_x2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      55.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END i0
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
        END
    END i4
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
        END
    END i5
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i3
    PIN i6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END i6
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 52.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 52.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 53.50 41.00 ;
    END
END oa3ao322_x2


MACRO oa3ao322_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      60.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END i2
    PIN i6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END i6
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
        END
    END i4
    PIN i5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
        END
    END i5
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i0
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 57.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 57.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 58.50 41.00 ;
    END
END oa3ao322_x4


MACRO on12_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
    END
END on12_x1


MACRO on12_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      40.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END q
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 37.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 37.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 38.50 41.00 ;
    END
END on12_x4


MACRO one_x0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      15.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END q
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 12.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 12.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 13.50 41.00 ;
    END
END one_x0


MACRO powmid_x0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 10.00 6.00 10.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 25.00 6.00 25.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
    END
END powmid_x0


MACRO rowend_x0
    CLASS     CORE FEEDTHRU ;
    ORIGIN    0.00 0.00 ;
    SIZE      5.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 2.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 2.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 3.50 41.00 ;
    END
END rowend_x0


MACRO sff1_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      90.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 79.00 39.00 81.00 41.00 ;
            RECT 79.00 34.00 81.00 36.00 ;
            RECT 79.00 29.00 81.00 31.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 79.00 19.00 81.00 21.00 ;
            RECT 79.00 14.00 81.00 16.00 ;
            RECT 79.00 9.00 81.00 11.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            LAYER L_ALU1 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END i
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END ck
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 87.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 87.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 88.50 41.00 ;
    END
END sff1_x4


MACRO sff2_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      120.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 109.00 39.00 111.00 41.00 ;
            RECT 109.00 34.00 111.00 36.00 ;
            RECT 109.00 29.00 111.00 31.00 ;
            RECT 109.00 24.00 111.00 26.00 ;
            RECT 109.00 19.00 111.00 21.00 ;
            RECT 109.00 14.00 111.00 16.00 ;
            RECT 109.00 9.00 111.00 11.00 ;
        END
    END q
    PIN cmd
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END cmd
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END i0
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
        END
    END ck
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 117.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 117.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 118.50 41.00 ;
    END
END sff2_x4


MACRO sff3_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      140.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 129.00 39.00 131.00 41.00 ;
            RECT 129.00 34.00 131.00 36.00 ;
            RECT 129.00 29.00 131.00 31.00 ;
            RECT 129.00 24.00 131.00 26.00 ;
            RECT 129.00 19.00 131.00 21.00 ;
            RECT 129.00 14.00 131.00 16.00 ;
            RECT 129.00 9.00 131.00 11.00 ;
        END
    END q
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END ck
    PIN cmd1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END cmd1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 24.00 26.00 26.00 ;
        END
    END i1
    PIN cmd0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END cmd0
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 19.00 41.00 21.00 ;
            LAYER L_ALU1 ;
            RECT 39.00 29.00 41.00 31.00 ;
            LAYER L_ALU1 ;
            RECT 44.00 24.00 46.00 26.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 137.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 137.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 138.50 41.00 ;
    END
END sff3_x4


MACRO tie_x0
    CLASS     CORE FEEDTHRU ;
    ORIGIN    0.00 0.00 ;
    SIZE      10.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 7.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 7.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 8.50 41.00 ;
    END
END tie_x0


MACRO ts_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END q
    PIN cmd
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END cmd
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
    END
END ts_x4


MACRO ts_x8
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      65.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU1 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 24.00 34.00 26.00 36.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 24.00 24.00 26.00 26.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 24.00 14.00 26.00 16.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END q
    PIN cmd
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
            RECT 29.00 9.00 31.00 11.00 ;
        END
    END cmd
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 54.00 34.00 56.00 36.00 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 54.00 24.00 56.00 26.00 ;
            RECT 54.00 19.00 56.00 21.00 ;
            RECT 54.00 14.00 56.00 16.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 62.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 62.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 63.50 41.00 ;
    END
END ts_x8


MACRO xr2_x1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 9.00 21.00 11.00 ;
            LAYER L_ALU1 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            LAYER L_ALU1 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 39.00 36.00 41.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
            RECT 34.00 9.00 36.00 11.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 43.50 41.00 ;
    END
END xr2_x1


MACRO xr2_x4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      60.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END q
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 34.00 39.00 36.00 41.00 ;
            RECT 34.00 34.00 36.00 36.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 34.00 24.00 36.00 26.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 57.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 57.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 58.50 41.00 ;
    END
END xr2_x4


MACRO zero_x0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      15.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 12.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 12.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 13.50 41.00 ;
    END
END zero_x0


END LIBRARY
