
MACRO rf2_dec_bufad0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END nq
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 29.00 26.00 31.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 43.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 43.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 43.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 43.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 43.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 43.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 43.50 41.00 ;
    END
END rf2_dec_bufad0


MACRO rf2_dec_bufad1_l
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END nq
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 31.00 21.00 ;
    END
END rf2_dec_bufad1_l


MACRO rf2_dec_bufad1_r
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      100.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END nq
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 97.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 97.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 51.00 11.00 ;
        RECT 54.00 9.00 56.00 11.00 ;
        RECT 59.00 9.00 61.00 11.00 ;
        RECT 64.00 9.00 66.00 11.00 ;
        RECT 69.00 9.00 71.00 11.00 ;
        RECT 74.00 9.00 76.00 11.00 ;
        RECT 79.00 9.00 81.00 11.00 ;
        RECT 84.00 9.00 86.00 11.00 ;
        RECT 89.00 9.00 91.00 11.00 ;
        RECT 94.00 9.00 98.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 51.00 16.00 ;
        RECT 54.00 14.00 56.00 16.00 ;
        RECT 59.00 14.00 61.00 16.00 ;
        RECT 64.00 14.00 66.00 16.00 ;
        RECT 69.00 14.00 71.00 16.00 ;
        RECT 74.00 14.00 76.00 16.00 ;
        RECT 79.00 14.00 81.00 16.00 ;
        RECT 84.00 14.00 86.00 16.00 ;
        RECT 89.00 14.00 91.00 16.00 ;
        RECT 94.00 14.00 98.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 51.00 21.00 ;
        RECT 54.00 19.00 56.00 21.00 ;
        RECT 59.00 19.00 61.00 21.00 ;
        RECT 64.00 19.00 66.00 21.00 ;
        RECT 69.00 19.00 71.00 21.00 ;
        RECT 74.00 19.00 76.00 21.00 ;
        RECT 79.00 19.00 81.00 21.00 ;
        RECT 84.00 19.00 86.00 21.00 ;
        RECT 89.00 19.00 91.00 21.00 ;
        RECT 94.00 19.00 98.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 51.00 26.00 ;
        RECT 54.00 24.00 56.00 26.00 ;
        RECT 59.00 24.00 61.00 26.00 ;
        RECT 64.00 24.00 66.00 26.00 ;
        RECT 69.00 24.00 71.00 26.00 ;
        RECT 74.00 24.00 76.00 26.00 ;
        RECT 79.00 24.00 81.00 26.00 ;
        RECT 84.00 24.00 86.00 26.00 ;
        RECT 89.00 24.00 91.00 26.00 ;
        RECT 94.00 24.00 98.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 51.00 31.00 ;
        RECT 54.00 29.00 56.00 31.00 ;
        RECT 59.00 29.00 61.00 31.00 ;
        RECT 64.00 29.00 66.00 31.00 ;
        RECT 69.00 29.00 71.00 31.00 ;
        RECT 74.00 29.00 76.00 31.00 ;
        RECT 79.00 29.00 81.00 31.00 ;
        RECT 84.00 29.00 86.00 31.00 ;
        RECT 89.00 29.00 91.00 31.00 ;
        RECT 94.00 29.00 98.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 51.00 36.00 ;
        RECT 54.00 34.00 56.00 36.00 ;
        RECT 59.00 34.00 61.00 36.00 ;
        RECT 64.00 34.00 66.00 36.00 ;
        RECT 69.00 34.00 71.00 36.00 ;
        RECT 74.00 34.00 76.00 36.00 ;
        RECT 79.00 34.00 81.00 36.00 ;
        RECT 84.00 34.00 86.00 36.00 ;
        RECT 89.00 34.00 91.00 36.00 ;
        RECT 94.00 34.00 98.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 51.00 41.00 ;
        RECT 54.00 39.00 56.00 41.00 ;
        RECT 59.00 39.00 61.00 41.00 ;
        RECT 64.00 39.00 66.00 41.00 ;
        RECT 69.00 39.00 71.00 41.00 ;
        RECT 74.00 39.00 76.00 41.00 ;
        RECT 79.00 39.00 81.00 41.00 ;
        RECT 84.00 39.00 86.00 41.00 ;
        RECT 89.00 39.00 91.00 41.00 ;
        RECT 94.00 39.00 98.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 31.00 21.00 ;
    END
END rf2_dec_bufad1_r


MACRO rf2_dec_bufad2_l
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq0
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END nq0
    PIN nq1
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END nq1
    PIN q0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END q0
    PIN q1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END q1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 48.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 48.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 48.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 48.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 48.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 48.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 48.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 46.00 21.00 ;
    END
END rf2_dec_bufad2_l


MACRO rf2_dec_bufad2_r
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      100.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq0
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END nq0
    PIN nq1
        DIRECTION INOUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END nq1
    PIN q0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END q0
    PIN q1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END q1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 97.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 97.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 51.00 11.00 ;
        RECT 54.00 9.00 56.00 11.00 ;
        RECT 59.00 9.00 61.00 11.00 ;
        RECT 64.00 9.00 66.00 11.00 ;
        RECT 69.00 9.00 71.00 11.00 ;
        RECT 74.00 9.00 76.00 11.00 ;
        RECT 79.00 9.00 81.00 11.00 ;
        RECT 84.00 9.00 86.00 11.00 ;
        RECT 89.00 9.00 91.00 11.00 ;
        RECT 94.00 9.00 98.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 51.00 16.00 ;
        RECT 54.00 14.00 56.00 16.00 ;
        RECT 59.00 14.00 61.00 16.00 ;
        RECT 64.00 14.00 66.00 16.00 ;
        RECT 69.00 14.00 71.00 16.00 ;
        RECT 74.00 14.00 76.00 16.00 ;
        RECT 79.00 14.00 81.00 16.00 ;
        RECT 84.00 14.00 86.00 16.00 ;
        RECT 89.00 14.00 91.00 16.00 ;
        RECT 94.00 14.00 98.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 51.00 21.00 ;
        RECT 54.00 19.00 56.00 21.00 ;
        RECT 59.00 19.00 61.00 21.00 ;
        RECT 64.00 19.00 66.00 21.00 ;
        RECT 69.00 19.00 71.00 21.00 ;
        RECT 74.00 19.00 76.00 21.00 ;
        RECT 79.00 19.00 81.00 21.00 ;
        RECT 84.00 19.00 86.00 21.00 ;
        RECT 89.00 19.00 91.00 21.00 ;
        RECT 94.00 19.00 98.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 51.00 26.00 ;
        RECT 54.00 24.00 56.00 26.00 ;
        RECT 59.00 24.00 61.00 26.00 ;
        RECT 64.00 24.00 66.00 26.00 ;
        RECT 69.00 24.00 71.00 26.00 ;
        RECT 74.00 24.00 76.00 26.00 ;
        RECT 79.00 24.00 81.00 26.00 ;
        RECT 84.00 24.00 86.00 26.00 ;
        RECT 89.00 24.00 91.00 26.00 ;
        RECT 94.00 24.00 98.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 51.00 31.00 ;
        RECT 54.00 29.00 56.00 31.00 ;
        RECT 59.00 29.00 61.00 31.00 ;
        RECT 64.00 29.00 66.00 31.00 ;
        RECT 69.00 29.00 71.00 31.00 ;
        RECT 74.00 29.00 76.00 31.00 ;
        RECT 79.00 29.00 81.00 31.00 ;
        RECT 84.00 29.00 86.00 31.00 ;
        RECT 89.00 29.00 91.00 31.00 ;
        RECT 94.00 29.00 98.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 51.00 36.00 ;
        RECT 54.00 34.00 56.00 36.00 ;
        RECT 59.00 34.00 61.00 36.00 ;
        RECT 64.00 34.00 66.00 36.00 ;
        RECT 69.00 34.00 71.00 36.00 ;
        RECT 74.00 34.00 76.00 36.00 ;
        RECT 79.00 34.00 81.00 36.00 ;
        RECT 84.00 34.00 86.00 36.00 ;
        RECT 89.00 34.00 91.00 36.00 ;
        RECT 94.00 34.00 98.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 51.00 41.00 ;
        RECT 54.00 39.00 56.00 41.00 ;
        RECT 59.00 39.00 61.00 41.00 ;
        RECT 64.00 39.00 66.00 41.00 ;
        RECT 69.00 39.00 71.00 41.00 ;
        RECT 74.00 39.00 76.00 41.00 ;
        RECT 79.00 39.00 81.00 41.00 ;
        RECT 84.00 39.00 86.00 41.00 ;
        RECT 89.00 39.00 91.00 41.00 ;
        RECT 94.00 39.00 98.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 46.00 21.00 ;
    END
END rf2_dec_bufad2_r


MACRO rf2_dec_nand2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      70.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 67.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 67.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 51.00 11.00 ;
        RECT 54.00 9.00 56.00 11.00 ;
        RECT 59.00 9.00 61.00 11.00 ;
        RECT 64.00 9.00 68.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 51.00 16.00 ;
        RECT 54.00 14.00 56.00 16.00 ;
        RECT 59.00 14.00 61.00 16.00 ;
        RECT 64.00 14.00 68.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 51.00 21.00 ;
        RECT 54.00 19.00 56.00 21.00 ;
        RECT 59.00 19.00 61.00 21.00 ;
        RECT 64.00 19.00 68.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 51.00 26.00 ;
        RECT 54.00 24.00 56.00 26.00 ;
        RECT 59.00 24.00 61.00 26.00 ;
        RECT 64.00 24.00 68.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 51.00 31.00 ;
        RECT 54.00 29.00 56.00 31.00 ;
        RECT 59.00 29.00 61.00 31.00 ;
        RECT 64.00 29.00 68.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 51.00 36.00 ;
        RECT 54.00 34.00 56.00 36.00 ;
        RECT 59.00 34.00 61.00 36.00 ;
        RECT 64.00 34.00 68.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 51.00 41.00 ;
        RECT 54.00 39.00 56.00 41.00 ;
        RECT 59.00 39.00 61.00 41.00 ;
        RECT 64.00 39.00 68.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 26.00 21.00 ;
        RECT 14.00 19.00 46.00 21.00 ;
    END
END rf2_dec_nand2


MACRO rf2_dec_nand3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      70.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 67.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 67.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 51.00 11.00 ;
        RECT 54.00 9.00 56.00 11.00 ;
        RECT 59.00 9.00 61.00 11.00 ;
        RECT 64.00 9.00 68.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 51.00 16.00 ;
        RECT 54.00 14.00 56.00 16.00 ;
        RECT 59.00 14.00 61.00 16.00 ;
        RECT 64.00 14.00 68.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 51.00 21.00 ;
        RECT 54.00 19.00 56.00 21.00 ;
        RECT 59.00 19.00 61.00 21.00 ;
        RECT 64.00 19.00 68.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 51.00 26.00 ;
        RECT 54.00 24.00 56.00 26.00 ;
        RECT 59.00 24.00 61.00 26.00 ;
        RECT 64.00 24.00 68.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 51.00 31.00 ;
        RECT 54.00 29.00 56.00 31.00 ;
        RECT 59.00 29.00 61.00 31.00 ;
        RECT 64.00 29.00 68.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 51.00 36.00 ;
        RECT 54.00 34.00 56.00 36.00 ;
        RECT 59.00 34.00 61.00 36.00 ;
        RECT 64.00 34.00 68.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 51.00 41.00 ;
        RECT 54.00 39.00 56.00 41.00 ;
        RECT 59.00 39.00 61.00 41.00 ;
        RECT 64.00 39.00 68.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 19.00 26.00 21.00 ;
        RECT 14.00 19.00 46.00 21.00 ;
    END
END rf2_dec_nand3


MACRO rf2_dec_nand4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      70.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END i2
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i0
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 67.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 67.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 51.00 11.00 ;
        RECT 54.00 9.00 56.00 11.00 ;
        RECT 59.00 9.00 61.00 11.00 ;
        RECT 64.00 9.00 68.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 51.00 16.00 ;
        RECT 54.00 14.00 56.00 16.00 ;
        RECT 59.00 14.00 61.00 16.00 ;
        RECT 64.00 14.00 68.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 51.00 21.00 ;
        RECT 54.00 19.00 56.00 21.00 ;
        RECT 59.00 19.00 61.00 21.00 ;
        RECT 64.00 19.00 68.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 51.00 26.00 ;
        RECT 54.00 24.00 56.00 26.00 ;
        RECT 59.00 24.00 61.00 26.00 ;
        RECT 64.00 24.00 68.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 51.00 31.00 ;
        RECT 54.00 29.00 56.00 31.00 ;
        RECT 59.00 29.00 61.00 31.00 ;
        RECT 64.00 29.00 68.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 51.00 36.00 ;
        RECT 54.00 34.00 56.00 36.00 ;
        RECT 59.00 34.00 61.00 36.00 ;
        RECT 64.00 34.00 68.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 51.00 41.00 ;
        RECT 54.00 39.00 56.00 41.00 ;
        RECT 59.00 39.00 61.00 41.00 ;
        RECT 64.00 39.00 68.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 14.00 19.00 46.00 21.00 ;
        RECT 19.00 19.00 26.00 21.00 ;
    END
END rf2_dec_nand4


MACRO rf2_dec_nao3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 39.00 11.00 41.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 34.00 21.00 36.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 33.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 33.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 33.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 33.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 33.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 33.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 33.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 19.00 11.00 21.00 ;
    END
END rf2_dec_nao3


MACRO rf2_dec_nbuf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      105.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 102.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 102.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 51.00 11.00 ;
        RECT 54.00 9.00 56.00 11.00 ;
        RECT 59.00 9.00 61.00 11.00 ;
        RECT 64.00 9.00 66.00 11.00 ;
        RECT 69.00 9.00 71.00 11.00 ;
        RECT 74.00 9.00 76.00 11.00 ;
        RECT 79.00 9.00 81.00 11.00 ;
        RECT 84.00 9.00 86.00 11.00 ;
        RECT 89.00 9.00 91.00 11.00 ;
        RECT 94.00 9.00 96.00 11.00 ;
        RECT 99.00 9.00 103.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 51.00 16.00 ;
        RECT 54.00 14.00 56.00 16.00 ;
        RECT 59.00 14.00 61.00 16.00 ;
        RECT 64.00 14.00 66.00 16.00 ;
        RECT 69.00 14.00 71.00 16.00 ;
        RECT 74.00 14.00 76.00 16.00 ;
        RECT 79.00 14.00 81.00 16.00 ;
        RECT 84.00 14.00 86.00 16.00 ;
        RECT 89.00 14.00 91.00 16.00 ;
        RECT 94.00 14.00 96.00 16.00 ;
        RECT 99.00 14.00 103.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 51.00 21.00 ;
        RECT 54.00 19.00 56.00 21.00 ;
        RECT 59.00 19.00 61.00 21.00 ;
        RECT 64.00 19.00 66.00 21.00 ;
        RECT 69.00 19.00 71.00 21.00 ;
        RECT 74.00 19.00 76.00 21.00 ;
        RECT 79.00 19.00 81.00 21.00 ;
        RECT 84.00 19.00 86.00 21.00 ;
        RECT 89.00 19.00 91.00 21.00 ;
        RECT 94.00 19.00 96.00 21.00 ;
        RECT 99.00 19.00 103.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 51.00 26.00 ;
        RECT 54.00 24.00 56.00 26.00 ;
        RECT 59.00 24.00 61.00 26.00 ;
        RECT 64.00 24.00 66.00 26.00 ;
        RECT 69.00 24.00 71.00 26.00 ;
        RECT 74.00 24.00 76.00 26.00 ;
        RECT 79.00 24.00 81.00 26.00 ;
        RECT 84.00 24.00 86.00 26.00 ;
        RECT 89.00 24.00 91.00 26.00 ;
        RECT 94.00 24.00 96.00 26.00 ;
        RECT 99.00 24.00 103.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 51.00 31.00 ;
        RECT 54.00 29.00 56.00 31.00 ;
        RECT 59.00 29.00 61.00 31.00 ;
        RECT 64.00 29.00 66.00 31.00 ;
        RECT 69.00 29.00 71.00 31.00 ;
        RECT 74.00 29.00 76.00 31.00 ;
        RECT 79.00 29.00 81.00 31.00 ;
        RECT 84.00 29.00 86.00 31.00 ;
        RECT 89.00 29.00 91.00 31.00 ;
        RECT 94.00 29.00 96.00 31.00 ;
        RECT 99.00 29.00 103.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 51.00 36.00 ;
        RECT 54.00 34.00 56.00 36.00 ;
        RECT 59.00 34.00 61.00 36.00 ;
        RECT 64.00 34.00 66.00 36.00 ;
        RECT 69.00 34.00 71.00 36.00 ;
        RECT 74.00 34.00 76.00 36.00 ;
        RECT 79.00 34.00 81.00 36.00 ;
        RECT 84.00 34.00 86.00 36.00 ;
        RECT 89.00 34.00 91.00 36.00 ;
        RECT 94.00 34.00 96.00 36.00 ;
        RECT 99.00 34.00 103.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 51.00 41.00 ;
        RECT 54.00 39.00 56.00 41.00 ;
        RECT 59.00 39.00 61.00 41.00 ;
        RECT 64.00 39.00 66.00 41.00 ;
        RECT 69.00 39.00 71.00 41.00 ;
        RECT 74.00 39.00 76.00 41.00 ;
        RECT 79.00 39.00 81.00 41.00 ;
        RECT 84.00 39.00 86.00 41.00 ;
        RECT 89.00 39.00 91.00 41.00 ;
        RECT 94.00 39.00 96.00 41.00 ;
        RECT 99.00 39.00 103.50 41.00 ;
    END
END rf2_dec_nbuf


MACRO rf2_dec_nor3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 39.00 11.00 41.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 33.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 33.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 33.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 33.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 33.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 33.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 33.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 19.00 11.00 21.00 ;
    END
END rf2_dec_nor3


MACRO rf2_inmux_buf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN sel0
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 39.00 36.00 41.00 ;
        END
    END sel0
    PIN sel1
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END sel1
    PIN sel
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 14.00 79.00 16.00 81.00 ;
            RECT 14.00 74.00 16.00 76.00 ;
            RECT 14.00 69.00 16.00 71.00 ;
        END
    END sel
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 42.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 42.00 97.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 43.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 43.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 43.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 43.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 43.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 43.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 43.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 21.00 61.00 ;
        RECT 24.00 59.00 26.00 61.00 ;
        RECT 29.00 59.00 31.00 61.00 ;
        RECT 34.00 59.00 36.00 61.00 ;
        RECT 39.00 59.00 43.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 26.00 66.00 ;
        RECT 29.00 64.00 31.00 66.00 ;
        RECT 34.00 64.00 36.00 66.00 ;
        RECT 39.00 64.00 43.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 21.00 71.00 ;
        RECT 24.00 69.00 26.00 71.00 ;
        RECT 29.00 69.00 31.00 71.00 ;
        RECT 34.00 69.00 36.00 71.00 ;
        RECT 39.00 69.00 43.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 21.00 76.00 ;
        RECT 24.00 74.00 26.00 76.00 ;
        RECT 29.00 74.00 31.00 76.00 ;
        RECT 34.00 74.00 36.00 76.00 ;
        RECT 39.00 74.00 43.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 21.00 81.00 ;
        RECT 24.00 79.00 26.00 81.00 ;
        RECT 29.00 79.00 31.00 81.00 ;
        RECT 34.00 79.00 36.00 81.00 ;
        RECT 39.00 79.00 43.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 21.00 86.00 ;
        RECT 24.00 84.00 26.00 86.00 ;
        RECT 29.00 84.00 31.00 86.00 ;
        RECT 34.00 84.00 36.00 86.00 ;
        RECT 39.00 84.00 43.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 21.00 91.00 ;
        RECT 24.00 89.00 26.00 91.00 ;
        RECT 29.00 89.00 31.00 91.00 ;
        RECT 34.00 89.00 36.00 91.00 ;
        RECT 39.00 89.00 43.50 91.00 ;
        LAYER L_ALU2 ;
        RECT 26.00 39.00 40.00 41.00 ;
        RECT 8.00 14.00 26.00 16.00 ;
        RECT 4.00 14.00 26.00 16.00 ;
        RECT 24.00 39.00 41.00 41.00 ;
    END
END rf2_inmux_buf


MACRO rf2_inmux_mem
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN dinx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END dinx
    PIN datain1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END datain1
    PIN datain0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END datain0
    PIN sel0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 29.00 36.00 31.00 ;
        END
    END sel0
    PIN sel1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 29.00 26.00 31.00 ;
        END
    END sel1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 43.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 43.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 43.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 43.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 43.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 43.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 43.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 24.00 29.00 36.00 31.00 ;
    END
END rf2_inmux_mem


MACRO rf2_mid_buf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN reada
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END reada
    PIN write
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END write
    PIN readb
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END readb
    PIN selrb
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 84.00 26.00 86.00 ;
        END
    END selrb
    PIN selra
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 84.00 16.00 86.00 ;
        END
    END selra
    PIN nck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT -1.00 89.00 1.00 91.00 ;
        END
    END nck
    PIN selw
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 84.00 11.00 86.00 ;
        END
    END selw
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 32.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 32.00 97.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 33.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 33.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 33.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 33.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 33.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 33.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 33.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 21.00 61.00 ;
        RECT 24.00 59.00 26.00 61.00 ;
        RECT 29.00 59.00 33.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 26.00 66.00 ;
        RECT 29.00 64.00 33.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 21.00 71.00 ;
        RECT 24.00 69.00 26.00 71.00 ;
        RECT 29.00 69.00 33.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 21.00 76.00 ;
        RECT 24.00 74.00 26.00 76.00 ;
        RECT 29.00 74.00 33.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 21.00 81.00 ;
        RECT 24.00 79.00 26.00 81.00 ;
        RECT 29.00 79.00 33.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 21.00 86.00 ;
        RECT 24.00 84.00 26.00 86.00 ;
        RECT 29.00 84.00 33.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 21.00 91.00 ;
        RECT 24.00 89.00 26.00 91.00 ;
        RECT 29.00 89.00 33.50 91.00 ;
        LAYER L_ALU2 ;
        RECT 14.00 64.00 31.00 66.00 ;
        RECT 4.00 59.00 31.00 61.00 ;
        RECT 4.00 39.00 31.00 41.00 ;
        RECT 14.00 19.00 26.00 21.00 ;
        RECT 4.00 14.00 31.00 16.00 ;
        RECT 17.00 39.00 21.00 41.00 ;
        RECT 17.00 14.00 21.00 16.00 ;
        RECT 14.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 31.00 66.00 ;
        LAYER L_ALU3 ;
        RECT 14.00 19.00 16.00 66.00 ;
        RECT 24.00 19.00 26.00 66.00 ;
        RECT 24.00 19.00 26.00 66.00 ;
        RECT 14.00 19.00 16.00 66.00 ;
    END
END rf2_mid_buf


MACRO rf2_mid_mem
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN busb
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 24.00 36.00 26.00 ;
        END
    END busb
    PIN busa
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END busa
    PIN write
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END write
    PIN dinx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END dinx
    PIN reada
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 29.00 21.00 31.00 ;
        END
    END reada
    PIN readb
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 29.00 31.00 31.00 ;
        END
    END readb
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 33.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 33.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 33.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 33.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 33.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 33.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 33.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 29.00 26.00 31.00 ;
        RECT 4.00 29.00 16.00 31.00 ;
    END
END rf2_mid_mem


MACRO rf2_mid_mem_r0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN busb
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 24.00 36.00 26.00 ;
        END
    END busb
    PIN busa
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER L_ALU2 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END busa
    PIN write
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END write
    PIN dinx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END dinx
    PIN reada
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 29.00 21.00 31.00 ;
        END
    END reada
    PIN readb
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 29.00 31.00 31.00 ;
        END
    END readb
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 33.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 33.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 33.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 33.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 33.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 33.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 33.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 19.00 29.00 26.00 31.00 ;
    END
END rf2_mid_mem_r0


MACRO rf2_out_buf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      105.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN xcks
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 59.00 16.00 61.00 ;
            RECT 14.00 54.00 16.00 56.00 ;
            RECT 14.00 49.00 16.00 51.00 ;
            RECT 14.00 44.00 16.00 46.00 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END xcks
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            LAYER L_ALU2 ;
            RECT 14.00 89.00 16.00 91.00 ;
        END
    END nck
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
        END
    END ck
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 102.00 47.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 102.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 102.00 3.00 ;
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 102.00 97.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 6.00 11.00 ;
        RECT 9.00 9.00 11.00 11.00 ;
        RECT 14.00 9.00 16.00 11.00 ;
        RECT 19.00 9.00 21.00 11.00 ;
        RECT 24.00 9.00 26.00 11.00 ;
        RECT 29.00 9.00 31.00 11.00 ;
        RECT 34.00 9.00 36.00 11.00 ;
        RECT 39.00 9.00 41.00 11.00 ;
        RECT 44.00 9.00 46.00 11.00 ;
        RECT 49.00 9.00 51.00 11.00 ;
        RECT 54.00 9.00 56.00 11.00 ;
        RECT 59.00 9.00 61.00 11.00 ;
        RECT 64.00 9.00 66.00 11.00 ;
        RECT 69.00 9.00 71.00 11.00 ;
        RECT 74.00 9.00 76.00 11.00 ;
        RECT 79.00 9.00 81.00 11.00 ;
        RECT 84.00 9.00 86.00 11.00 ;
        RECT 89.00 9.00 91.00 11.00 ;
        RECT 94.00 9.00 96.00 11.00 ;
        RECT 99.00 9.00 103.50 11.00 ;
        RECT 1.50 14.00 6.00 16.00 ;
        RECT 9.00 14.00 11.00 16.00 ;
        RECT 14.00 14.00 16.00 16.00 ;
        RECT 19.00 14.00 21.00 16.00 ;
        RECT 24.00 14.00 26.00 16.00 ;
        RECT 29.00 14.00 31.00 16.00 ;
        RECT 34.00 14.00 36.00 16.00 ;
        RECT 39.00 14.00 41.00 16.00 ;
        RECT 44.00 14.00 46.00 16.00 ;
        RECT 49.00 14.00 51.00 16.00 ;
        RECT 54.00 14.00 56.00 16.00 ;
        RECT 59.00 14.00 61.00 16.00 ;
        RECT 64.00 14.00 66.00 16.00 ;
        RECT 69.00 14.00 71.00 16.00 ;
        RECT 74.00 14.00 76.00 16.00 ;
        RECT 79.00 14.00 81.00 16.00 ;
        RECT 84.00 14.00 86.00 16.00 ;
        RECT 89.00 14.00 91.00 16.00 ;
        RECT 94.00 14.00 96.00 16.00 ;
        RECT 99.00 14.00 103.50 16.00 ;
        RECT 1.50 19.00 6.00 21.00 ;
        RECT 9.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 16.00 21.00 ;
        RECT 19.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 26.00 21.00 ;
        RECT 29.00 19.00 31.00 21.00 ;
        RECT 34.00 19.00 36.00 21.00 ;
        RECT 39.00 19.00 41.00 21.00 ;
        RECT 44.00 19.00 46.00 21.00 ;
        RECT 49.00 19.00 51.00 21.00 ;
        RECT 54.00 19.00 56.00 21.00 ;
        RECT 59.00 19.00 61.00 21.00 ;
        RECT 64.00 19.00 66.00 21.00 ;
        RECT 69.00 19.00 71.00 21.00 ;
        RECT 74.00 19.00 76.00 21.00 ;
        RECT 79.00 19.00 81.00 21.00 ;
        RECT 84.00 19.00 86.00 21.00 ;
        RECT 89.00 19.00 91.00 21.00 ;
        RECT 94.00 19.00 96.00 21.00 ;
        RECT 99.00 19.00 103.50 21.00 ;
        RECT 1.50 24.00 6.00 26.00 ;
        RECT 9.00 24.00 11.00 26.00 ;
        RECT 14.00 24.00 16.00 26.00 ;
        RECT 19.00 24.00 21.00 26.00 ;
        RECT 24.00 24.00 26.00 26.00 ;
        RECT 29.00 24.00 31.00 26.00 ;
        RECT 34.00 24.00 36.00 26.00 ;
        RECT 39.00 24.00 41.00 26.00 ;
        RECT 44.00 24.00 46.00 26.00 ;
        RECT 49.00 24.00 51.00 26.00 ;
        RECT 54.00 24.00 56.00 26.00 ;
        RECT 59.00 24.00 61.00 26.00 ;
        RECT 64.00 24.00 66.00 26.00 ;
        RECT 69.00 24.00 71.00 26.00 ;
        RECT 74.00 24.00 76.00 26.00 ;
        RECT 79.00 24.00 81.00 26.00 ;
        RECT 84.00 24.00 86.00 26.00 ;
        RECT 89.00 24.00 91.00 26.00 ;
        RECT 94.00 24.00 96.00 26.00 ;
        RECT 99.00 24.00 103.50 26.00 ;
        RECT 1.50 29.00 6.00 31.00 ;
        RECT 9.00 29.00 11.00 31.00 ;
        RECT 14.00 29.00 16.00 31.00 ;
        RECT 19.00 29.00 21.00 31.00 ;
        RECT 24.00 29.00 26.00 31.00 ;
        RECT 29.00 29.00 31.00 31.00 ;
        RECT 34.00 29.00 36.00 31.00 ;
        RECT 39.00 29.00 41.00 31.00 ;
        RECT 44.00 29.00 46.00 31.00 ;
        RECT 49.00 29.00 51.00 31.00 ;
        RECT 54.00 29.00 56.00 31.00 ;
        RECT 59.00 29.00 61.00 31.00 ;
        RECT 64.00 29.00 66.00 31.00 ;
        RECT 69.00 29.00 71.00 31.00 ;
        RECT 74.00 29.00 76.00 31.00 ;
        RECT 79.00 29.00 81.00 31.00 ;
        RECT 84.00 29.00 86.00 31.00 ;
        RECT 89.00 29.00 91.00 31.00 ;
        RECT 94.00 29.00 96.00 31.00 ;
        RECT 99.00 29.00 103.50 31.00 ;
        RECT 1.50 34.00 6.00 36.00 ;
        RECT 9.00 34.00 11.00 36.00 ;
        RECT 14.00 34.00 16.00 36.00 ;
        RECT 19.00 34.00 21.00 36.00 ;
        RECT 24.00 34.00 26.00 36.00 ;
        RECT 29.00 34.00 31.00 36.00 ;
        RECT 34.00 34.00 36.00 36.00 ;
        RECT 39.00 34.00 41.00 36.00 ;
        RECT 44.00 34.00 46.00 36.00 ;
        RECT 49.00 34.00 51.00 36.00 ;
        RECT 54.00 34.00 56.00 36.00 ;
        RECT 59.00 34.00 61.00 36.00 ;
        RECT 64.00 34.00 66.00 36.00 ;
        RECT 69.00 34.00 71.00 36.00 ;
        RECT 74.00 34.00 76.00 36.00 ;
        RECT 79.00 34.00 81.00 36.00 ;
        RECT 84.00 34.00 86.00 36.00 ;
        RECT 89.00 34.00 91.00 36.00 ;
        RECT 94.00 34.00 96.00 36.00 ;
        RECT 99.00 34.00 103.50 36.00 ;
        RECT 1.50 39.00 6.00 41.00 ;
        RECT 9.00 39.00 11.00 41.00 ;
        RECT 14.00 39.00 16.00 41.00 ;
        RECT 19.00 39.00 21.00 41.00 ;
        RECT 24.00 39.00 26.00 41.00 ;
        RECT 29.00 39.00 31.00 41.00 ;
        RECT 34.00 39.00 36.00 41.00 ;
        RECT 39.00 39.00 41.00 41.00 ;
        RECT 44.00 39.00 46.00 41.00 ;
        RECT 49.00 39.00 51.00 41.00 ;
        RECT 54.00 39.00 56.00 41.00 ;
        RECT 59.00 39.00 61.00 41.00 ;
        RECT 64.00 39.00 66.00 41.00 ;
        RECT 69.00 39.00 71.00 41.00 ;
        RECT 74.00 39.00 76.00 41.00 ;
        RECT 79.00 39.00 81.00 41.00 ;
        RECT 84.00 39.00 86.00 41.00 ;
        RECT 89.00 39.00 91.00 41.00 ;
        RECT 94.00 39.00 96.00 41.00 ;
        RECT 99.00 39.00 103.50 41.00 ;
        RECT 1.50 59.00 6.00 61.00 ;
        RECT 9.00 59.00 11.00 61.00 ;
        RECT 14.00 59.00 16.00 61.00 ;
        RECT 19.00 59.00 21.00 61.00 ;
        RECT 24.00 59.00 26.00 61.00 ;
        RECT 29.00 59.00 31.00 61.00 ;
        RECT 34.00 59.00 36.00 61.00 ;
        RECT 39.00 59.00 41.00 61.00 ;
        RECT 44.00 59.00 46.00 61.00 ;
        RECT 49.00 59.00 51.00 61.00 ;
        RECT 54.00 59.00 56.00 61.00 ;
        RECT 59.00 59.00 61.00 61.00 ;
        RECT 64.00 59.00 66.00 61.00 ;
        RECT 69.00 59.00 71.00 61.00 ;
        RECT 74.00 59.00 76.00 61.00 ;
        RECT 79.00 59.00 81.00 61.00 ;
        RECT 84.00 59.00 86.00 61.00 ;
        RECT 89.00 59.00 91.00 61.00 ;
        RECT 94.00 59.00 96.00 61.00 ;
        RECT 99.00 59.00 103.50 61.00 ;
        RECT 1.50 64.00 6.00 66.00 ;
        RECT 9.00 64.00 11.00 66.00 ;
        RECT 14.00 64.00 16.00 66.00 ;
        RECT 19.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 26.00 66.00 ;
        RECT 29.00 64.00 31.00 66.00 ;
        RECT 34.00 64.00 36.00 66.00 ;
        RECT 39.00 64.00 41.00 66.00 ;
        RECT 44.00 64.00 46.00 66.00 ;
        RECT 49.00 64.00 51.00 66.00 ;
        RECT 54.00 64.00 56.00 66.00 ;
        RECT 59.00 64.00 61.00 66.00 ;
        RECT 64.00 64.00 66.00 66.00 ;
        RECT 69.00 64.00 71.00 66.00 ;
        RECT 74.00 64.00 76.00 66.00 ;
        RECT 79.00 64.00 81.00 66.00 ;
        RECT 84.00 64.00 86.00 66.00 ;
        RECT 89.00 64.00 91.00 66.00 ;
        RECT 94.00 64.00 96.00 66.00 ;
        RECT 99.00 64.00 103.50 66.00 ;
        RECT 1.50 69.00 6.00 71.00 ;
        RECT 9.00 69.00 11.00 71.00 ;
        RECT 14.00 69.00 16.00 71.00 ;
        RECT 19.00 69.00 21.00 71.00 ;
        RECT 24.00 69.00 26.00 71.00 ;
        RECT 29.00 69.00 31.00 71.00 ;
        RECT 34.00 69.00 36.00 71.00 ;
        RECT 39.00 69.00 41.00 71.00 ;
        RECT 44.00 69.00 46.00 71.00 ;
        RECT 49.00 69.00 51.00 71.00 ;
        RECT 54.00 69.00 56.00 71.00 ;
        RECT 59.00 69.00 61.00 71.00 ;
        RECT 64.00 69.00 66.00 71.00 ;
        RECT 69.00 69.00 71.00 71.00 ;
        RECT 74.00 69.00 76.00 71.00 ;
        RECT 79.00 69.00 81.00 71.00 ;
        RECT 84.00 69.00 86.00 71.00 ;
        RECT 89.00 69.00 91.00 71.00 ;
        RECT 94.00 69.00 96.00 71.00 ;
        RECT 99.00 69.00 103.50 71.00 ;
        RECT 1.50 74.00 6.00 76.00 ;
        RECT 9.00 74.00 11.00 76.00 ;
        RECT 14.00 74.00 16.00 76.00 ;
        RECT 19.00 74.00 21.00 76.00 ;
        RECT 24.00 74.00 26.00 76.00 ;
        RECT 29.00 74.00 31.00 76.00 ;
        RECT 34.00 74.00 36.00 76.00 ;
        RECT 39.00 74.00 41.00 76.00 ;
        RECT 44.00 74.00 46.00 76.00 ;
        RECT 49.00 74.00 51.00 76.00 ;
        RECT 54.00 74.00 56.00 76.00 ;
        RECT 59.00 74.00 61.00 76.00 ;
        RECT 64.00 74.00 66.00 76.00 ;
        RECT 69.00 74.00 71.00 76.00 ;
        RECT 74.00 74.00 76.00 76.00 ;
        RECT 79.00 74.00 81.00 76.00 ;
        RECT 84.00 74.00 86.00 76.00 ;
        RECT 89.00 74.00 91.00 76.00 ;
        RECT 94.00 74.00 96.00 76.00 ;
        RECT 99.00 74.00 103.50 76.00 ;
        RECT 1.50 79.00 6.00 81.00 ;
        RECT 9.00 79.00 11.00 81.00 ;
        RECT 14.00 79.00 16.00 81.00 ;
        RECT 19.00 79.00 21.00 81.00 ;
        RECT 24.00 79.00 26.00 81.00 ;
        RECT 29.00 79.00 31.00 81.00 ;
        RECT 34.00 79.00 36.00 81.00 ;
        RECT 39.00 79.00 41.00 81.00 ;
        RECT 44.00 79.00 46.00 81.00 ;
        RECT 49.00 79.00 51.00 81.00 ;
        RECT 54.00 79.00 56.00 81.00 ;
        RECT 59.00 79.00 61.00 81.00 ;
        RECT 64.00 79.00 66.00 81.00 ;
        RECT 69.00 79.00 71.00 81.00 ;
        RECT 74.00 79.00 76.00 81.00 ;
        RECT 79.00 79.00 81.00 81.00 ;
        RECT 84.00 79.00 86.00 81.00 ;
        RECT 89.00 79.00 91.00 81.00 ;
        RECT 94.00 79.00 96.00 81.00 ;
        RECT 99.00 79.00 103.50 81.00 ;
        RECT 1.50 84.00 6.00 86.00 ;
        RECT 9.00 84.00 11.00 86.00 ;
        RECT 14.00 84.00 16.00 86.00 ;
        RECT 19.00 84.00 21.00 86.00 ;
        RECT 24.00 84.00 26.00 86.00 ;
        RECT 29.00 84.00 31.00 86.00 ;
        RECT 34.00 84.00 36.00 86.00 ;
        RECT 39.00 84.00 41.00 86.00 ;
        RECT 44.00 84.00 46.00 86.00 ;
        RECT 49.00 84.00 51.00 86.00 ;
        RECT 54.00 84.00 56.00 86.00 ;
        RECT 59.00 84.00 61.00 86.00 ;
        RECT 64.00 84.00 66.00 86.00 ;
        RECT 69.00 84.00 71.00 86.00 ;
        RECT 74.00 84.00 76.00 86.00 ;
        RECT 79.00 84.00 81.00 86.00 ;
        RECT 84.00 84.00 86.00 86.00 ;
        RECT 89.00 84.00 91.00 86.00 ;
        RECT 94.00 84.00 96.00 86.00 ;
        RECT 99.00 84.00 103.50 86.00 ;
        RECT 1.50 89.00 6.00 91.00 ;
        RECT 9.00 89.00 11.00 91.00 ;
        RECT 14.00 89.00 16.00 91.00 ;
        RECT 19.00 89.00 21.00 91.00 ;
        RECT 24.00 89.00 26.00 91.00 ;
        RECT 29.00 89.00 31.00 91.00 ;
        RECT 34.00 89.00 36.00 91.00 ;
        RECT 39.00 89.00 41.00 91.00 ;
        RECT 44.00 89.00 46.00 91.00 ;
        RECT 49.00 89.00 51.00 91.00 ;
        RECT 54.00 89.00 56.00 91.00 ;
        RECT 59.00 89.00 61.00 91.00 ;
        RECT 64.00 89.00 66.00 91.00 ;
        RECT 69.00 89.00 71.00 91.00 ;
        RECT 74.00 89.00 76.00 91.00 ;
        RECT 79.00 89.00 81.00 91.00 ;
        RECT 84.00 89.00 86.00 91.00 ;
        RECT 89.00 89.00 91.00 91.00 ;
        RECT 94.00 89.00 96.00 91.00 ;
        RECT 99.00 89.00 103.50 91.00 ;
        LAYER L_ALU2 ;
        RECT 9.00 59.00 21.00 61.00 ;
        RECT 9.00 39.00 21.00 41.00 ;
        RECT 9.00 14.00 21.00 16.00 ;
    END
END rf2_out_buf

