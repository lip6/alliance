#
# $Id: cmos.lef,v 1.5 2004/09/29 21:40:39 jpc Exp $
#
# /------------------------------------------------------------------\
# |                                                                  |
# |        A l l i a n c e   C A D   S y s t e m                     |
# |  S i l i c o n   E n s e m b l e / A l l i a n c e               |
# |                                                                  |
# |  Author    :                      Jean-Paul CHAPUT               |
# |  E-mail    :         alliance-users@asim.lip6.fr                 |
# | ================================================================ |
# |  LEF       :         "./cmos_12.lef"                             |
# | **************************************************************** |
# |  U p d a t e s                                                   |
# |                                                                  |
# \------------------------------------------------------------------/
#


VERSION               5.2 ;
NAMESCASESENSITIVE    ON ;
BUSBITCHARS           "()" ;
DIVIDERCHAR           "." ;

#NOWIREEXTENSIONATPIN ON ;


UNITS
    DATABASE MICRONS 100  ;
END UNITS


LAYER POLY
    TYPE MASTERSLICE ;
END POLY


LAYER VIAP
    TYPE CUT ;
END VIAP


LAYER ALU1
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END ALU1


LAYER VIA1
    TYPE CUT ;
END VIA1


LAYER ALU2
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END ALU2


LAYER VIA2
    TYPE CUT ;
END VIA2


LAYER ALU3
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END ALU3


LAYER VIA3
    TYPE CUT ;
END VIA3


LAYER ALU4
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END ALU4


LAYER VIA4
    TYPE CUT ;
END VIA4


LAYER ALU5
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END ALU5


LAYER VIA5
    TYPE CUT ;
END VIA5


LAYER ALU6
    TYPE ROUTING ;
    WIDTH 2.00 ;
    SPACING 3.00 ;
    PITCH 5.00 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000032 ;
    RESISTANCE RPERSQ 0.100000 ;
END ALU6


#VIA CONT_POLY DEFAULT
#    LAYER POLY ;
#        RECT -1.50 -1.50 1.50 1.50 ;
#    LAYER VIAP ;
#        RECT -0.50 -0.50 0.50 0.50 ;
#    LAYER ALU1 ;
#        RECT -1.00 -1.00 1.00 1.00 ;
#END CONT_POLY


VIA CONT_VIA DEFAULT
    LAYER ALU1 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER VIA1 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER ALU2 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA


VIA CONT_VIA2 DEFAULT
    LAYER ALU3 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER VIA2 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER ALU2 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA2


VIA CONT_VIA3 DEFAULT
    LAYER ALU4 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER VIA3 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER ALU3 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA3


VIA CONT_VIA4 DEFAULT
    LAYER ALU5 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER VIA4 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER ALU4 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA4


VIA CONT_VIA5 DEFAULT
    LAYER ALU6 ;
        RECT -1.00 -1.00 1.00 1.00 ;
    LAYER VIA5 ;
        RECT -0.50 -0.50 0.50 0.50 ;
    LAYER ALU5 ;
        RECT -1.00 -1.00 1.00 1.00 ;
END CONT_VIA5


VIARULE TURN_ALU1 GENERATE
    LAYER ALU1 ;
        DIRECTION vertical ;

    LAYER ALU1 ;
        DIRECTION horizontal ;
END TURN_ALU1


VIARULE TURN_ALU2 GENERATE
    LAYER ALU2 ;
        DIRECTION vertical ;

    LAYER ALU2 ;
        DIRECTION horizontal ;
END TURN_ALU2


VIARULE TURN_ALU3 GENERATE
    LAYER ALU3 ;
        DIRECTION vertical ;

    LAYER ALU3 ;
        DIRECTION horizontal ;
END TURN_ALU3


VIARULE TURN_ALU4 GENERATE
    LAYER ALU4 ;
        DIRECTION vertical ;

    LAYER ALU4 ;
        DIRECTION horizontal ;
END TURN_ALU4


VIARULE TURN_ALU5 GENERATE
    LAYER ALU5 ;
        DIRECTION vertical ;

    LAYER ALU5 ;
        DIRECTION horizontal ;
END TURN_ALU5


VIARULE TURN_ALU6 GENERATE
    LAYER ALU6 ;
        DIRECTION vertical ;

    LAYER ALU6 ;
        DIRECTION horizontal ;
END TURN_ALU6


#VIARULE VIA1_HV
#    LAYER ALU1 ;
#        DIRECTION VERTICAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    LAYER ALU2 ;
#        DIRECTION HORIZONTAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    VIA CONT_VIA ;
#END VIA1_HV
#
#
#VIARULE VIA2_VH
#    LAYER ALU2 ;
#        DIRECTION HORIZONTAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    LAYER ALU3 ;
#        DIRECTION VERTICAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    VIA CONT_VIA2 ;
#END VIA2_VH
#
#
#VIARULE VIA3_VH
#    LAYER ALU3 ;
#        DIRECTION HORIZONTAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    LAYER ALU4 ;
#        DIRECTION VERTICAL ;
#        OVERHANG 0.50 ;
#        METALOVERHANG 0.50 ;
#
#    VIA CONT_VIA3 ;
#END VIA3_VH


VIARULE genVIA1_HV GENERATE
    LAYER ALU1 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER ALU2 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER VIA1 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA1_HV


VIARULE genVIA1_VH GENERATE
    LAYER ALU1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER ALU2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER VIA1 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA1_VH


VIARULE genVIA2_VH GENERATE
    LAYER ALU2 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER ALU3 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER VIA2 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA2_VH


VIARULE genVIA2_HV GENERATE
    LAYER ALU2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER ALU3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER VIA2 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA2_HV


VIARULE genVIA3_VH GENERATE
    LAYER ALU3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER ALU4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER VIA3 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA3_VH


VIARULE genVIA3_HV GENERATE
    LAYER ALU3 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER ALU4 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.50 ;
        METALOVERHANG 0.50 ;

    LAYER VIA3 ;
        RECT -0.50 -0.50 0.50 0.50 ;
        SPACING 3.00 BY 3.00 ;
END genVIA3_HV


SPACING
    SAMENET VIAP VIAP 3.00 ;
    SAMENET VIA1 VIA1 3.00 ;
    SAMENET VIA2 VIA2 3.00 ;
    SAMENET VIAP VIA1 3.00 STACK ;
    SAMENET VIA1 VIA2 3.00 STACK ;
    SAMENET VIA2 VIA3 3.00 STACK ;
    SAMENET VIA3 VIA4 3.00 STACK ;
    SAMENET VIA4 VIA5 3.00 STACK ;
    SAMENET POLY POLY 3.00 ;
    SAMENET ALU1 ALU1 3.00 STACK ;
    SAMENET ALU2 ALU2 3.00 STACK ;
    SAMENET ALU3 ALU3 3.00 STACK ;
    SAMENET ALU4 ALU4 3.00 STACK ;
    SAMENET ALU5 ALU5 3.00 STACK ;
    SAMENET ALU6 ALU6 3.00 ;
END SPACING


SITE core
    SYMMETRY y  ;
    CLASS CORE  ;
    SIZE 5.00 BY 50.00 ;
END core


SITE pad
    SYMMETRY y  ;
    CLASS PAD  ;
    SIZE 1.00 BY 500.00 ;
END pad


SITE corner
    SYMMETRY y r90  ;
    CLASS PAD  ;
    SIZE 500.00 BY 500.00 ;
END corner


END LIBRARY
