
MACRO ram_mem_buf0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 0.00 6.00 0.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 25.00 6.00 25.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 10.00 24.00 16.00 26.00 ;
        RECT 5.00 19.00 19.00 21.00 ;
        RECT 10.00 24.00 16.00 26.00 ;
        RECT 5.00 19.00 19.00 21.00 ;
    END
END ram_mem_buf0


MACRO ram_mem_buf1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nseli
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 34.00 16.00 36.00 ;
        END
    END nseli
    PIN nck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 9.00 24.00 11.00 26.00 ;
        END
    END nck
    PIN selramx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
        END
    END selramx
    PIN seli
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END seli
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 0.00 6.00 0.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 25.00 6.00 25.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 9.00 14.00 16.00 16.00 ;
        RECT 9.00 14.00 16.00 16.00 ;
        RECT 9.00 34.00 16.00 36.00 ;
        RECT 9.00 34.00 16.00 36.00 ;
    END
END ram_mem_buf1


MACRO ram_mem_data
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN selxi
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 44.00 11.00 46.00 ;
        END
    END selxi
    PIN bit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
            RECT -1.00 9.00 1.00 11.00 ;
        END
    END bit0
    PIN nbit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 19.00 26.00 21.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT -1.00 19.00 1.00 21.00 ;
        END
    END nbit0
    PIN nbit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT -1.00 39.00 1.00 41.00 ;
        END
    END nbit1
    PIN bit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT -1.00 29.00 1.00 31.00 ;
        END
    END bit1
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 25.00 6.00 25.00 44.00 ;
        END
    END vss
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 0.00 6.00 0.00 44.00 ;
        END
    END vdd
    OBS
        LAYER L_ALU2 ;
        RECT 24.00 37.00 26.00 41.00 ;
        RECT 24.00 29.00 26.00 33.00 ;
        RECT 24.00 9.00 26.00 15.00 ;
        RECT -1.00 4.00 26.00 46.00 ;
        RECT 19.00 4.00 26.00 6.00 ;
        RECT 19.00 24.00 26.00 26.00 ;
        RECT -1.00 24.00 6.00 26.00 ;
        RECT -1.00 14.00 6.00 16.00 ;
        RECT 19.00 44.00 26.00 46.00 ;
        RECT 9.00 44.00 16.00 46.00 ;
    END
END ram_mem_data


MACRO ram_mem_dec2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      100.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN ndeca
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END ndeca
    PIN ndecb
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 19.00 86.00 21.00 ;
        END
    END ndecb
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 19.00 61.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 97.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 25.00 6.00 25.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 75.00 6.00 75.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 97.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 0.00 6.00 0.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 50.00 6.00 50.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 100.00 6.00 100.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 98.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 29.00 19.00 36.00 21.00 ;
        RECT 79.00 19.00 86.00 21.00 ;
        RECT 59.00 19.00 66.00 21.00 ;
        RECT 9.00 19.00 16.00 21.00 ;
        RECT 9.00 19.00 86.00 21.00 ;
    END
END ram_mem_dec2


MACRO ram_mem_dec3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      100.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN ndeca
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END ndeca
    PIN ndecb
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 19.00 86.00 21.00 ;
        END
    END ndecb
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 19.00 61.00 21.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 97.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 25.00 6.00 25.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 75.00 6.00 75.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 97.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 0.00 6.00 0.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 50.00 6.00 50.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 100.00 6.00 100.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 98.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 19.00 11.00 21.00 ;
        RECT 14.00 19.00 21.00 21.00 ;
        RECT 29.00 19.00 36.00 21.00 ;
        RECT 54.00 19.00 61.00 21.00 ;
        RECT 79.00 19.00 86.00 21.00 ;
        RECT 4.00 19.00 86.00 21.00 ;
    END
END ram_mem_dec3


MACRO ram_mem_dec4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      100.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN ndeca
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END ndeca
    PIN ndecb
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 19.00 86.00 21.00 ;
        END
    END ndecb
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 19.00 66.00 21.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 19.00 61.00 21.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 97.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 25.00 6.00 25.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 75.00 6.00 75.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 97.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 0.00 6.00 0.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 50.00 6.00 50.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 100.00 6.00 100.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 98.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 79.00 19.00 86.00 21.00 ;
        RECT 64.00 19.00 71.00 21.00 ;
        RECT 54.00 19.00 61.00 21.00 ;
        RECT 29.00 19.00 36.00 21.00 ;
        RECT 14.00 19.00 21.00 21.00 ;
        RECT 4.00 19.00 11.00 21.00 ;
        RECT 4.00 19.00 86.00 21.00 ;
    END
END ram_mem_dec4


MACRO ram_mem_dec5
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      100.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN ndecb
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 84.00 19.00 86.00 21.00 ;
        END
    END ndecb
    PIN ndeca
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END ndeca
    PIN i4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 19.00 66.00 21.00 ;
        END
    END i4
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 59.00 19.00 61.00 21.00 ;
        END
    END i3
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 9.00 19.00 11.00 21.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 97.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 25.00 6.00 25.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 75.00 6.00 75.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 97.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 0.00 6.00 0.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 50.00 6.00 50.00 44.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 100.00 6.00 100.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 98.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 79.00 19.00 86.00 21.00 ;
        RECT 64.00 19.00 71.00 21.00 ;
        RECT 54.00 19.00 61.00 21.00 ;
        RECT 39.00 19.00 46.00 21.00 ;
        RECT 29.00 19.00 36.00 21.00 ;
        RECT 4.00 19.00 86.00 21.00 ;
        RECT 14.00 19.00 21.00 21.00 ;
        RECT 4.00 19.00 11.00 21.00 ;
    END
END ram_mem_dec5


MACRO ram_mem_deci
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      25.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN seli
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 9.00 16.00 11.00 ;
        END
    END seli
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 9.00 34.00 11.00 36.00 ;
        END
    END i0
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 22.00 47.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 0.00 6.00 0.00 44.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 22.00 3.00 ;
            LAYER L_ALU3 ;
            WIDTH 12.00 ;
            PATH 25.00 6.00 25.00 44.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 23.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 9.00 9.00 16.00 11.00 ;
        RECT 9.00 9.00 16.00 11.00 ;
    END
END ram_mem_deci


MACRO ram_prech_buf0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 24.00 21.00 26.00 ;
        END
    END i
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 14.00 19.00 21.00 21.00 ;
        RECT 14.00 24.00 21.00 26.00 ;
        RECT 14.00 24.00 21.00 26.00 ;
        RECT 14.00 19.00 21.00 21.00 ;
        LAYER L_ALU3 ;
        RECT 4.00 -1.00 16.00 51.00 ;
        RECT 24.00 -1.00 36.00 51.00 ;
    END
END ram_prech_buf0


MACRO ram_prech_buf1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nckx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 34.00 21.00 36.00 ;
        END
    END nckx
    PIN nck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END nck
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 9.00 34.00 21.00 36.00 ;
        RECT 9.00 34.00 21.00 36.00 ;
        RECT 4.00 44.00 31.00 56.00 ;
        RECT 4.00 -6.00 31.00 6.00 ;
        LAYER L_ALU3 ;
        RECT 24.00 -1.00 36.00 51.00 ;
        RECT 4.00 -1.00 16.00 51.00 ;
    END
END ram_prech_buf1


MACRO ram_prech_data
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nbit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END nbit0
    PIN nbit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 24.00 39.00 26.00 41.00 ;
        END
    END nbit1
    PIN bit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
        END
    END bit1
    PIN bit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 29.00 9.00 31.00 11.00 ;
            RECT 24.00 9.00 26.00 11.00 ;
        END
    END bit0
    PIN prech
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END prech
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE FEEDTHRU ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 7.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE FEEDTHRU ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 7.00 3.00 ;
            PATH 23.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 13.00 0.00 17.00 6.00 ;
        RECT 1.50 9.00 28.50 41.00 ;
        RECT 13.00 44.00 28.50 50.00 ;
        LAYER L_ALU2 ;
        RECT 4.00 9.00 21.00 41.00 ;
        RECT 4.00 39.00 21.00 41.00 ;
        RECT 4.00 21.00 21.00 23.00 ;
        RECT 4.00 15.00 21.00 17.00 ;
        RECT 4.00 33.00 21.00 35.00 ;
        RECT 9.00 27.00 15.00 29.00 ;
        RECT 9.00 9.00 15.00 11.00 ;
        LAYER L_ALU3 ;
        RECT 4.00 -1.00 16.00 51.00 ;
        RECT 24.00 -1.00 36.00 51.00 ;
    END
END ram_prech_data


MACRO ram_prech_dec0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      30.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 27.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 27.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 28.50 41.00 ;
        LAYER L_ALU3 ;
        RECT 4.00 -1.00 16.00 51.00 ;
        RECT 24.00 -1.00 36.00 51.00 ;
    END
END ram_prech_dec0


MACRO ram_sense_buf0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      170.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN prech
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 19.00 116.00 21.00 ;
        END
    END prech
    PIN nsensex
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 24.00 91.00 26.00 ;
        END
    END nsensex
    PIN writex
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 134.00 24.00 136.00 26.00 ;
        END
    END writex
    PIN sensex
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 74.00 19.00 76.00 21.00 ;
        END
    END sensex
    PIN nad0x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END nad0x
    PIN ad0x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 24.00 31.00 26.00 ;
        END
    END ad0x
    PIN nckx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 104.00 24.00 106.00 26.00 ;
        END
    END nckx
    PIN ad0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END ad0
    PIN nwrite
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 139.00 19.00 141.00 21.00 ;
        END
    END nwrite
    PIN nsense
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 24.00 71.00 26.00 ;
        END
    END nsense
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 167.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 167.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 168.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 14.00 19.00 141.00 21.00 ;
        RECT 64.00 24.00 71.00 26.00 ;
        RECT 104.00 24.00 111.00 26.00 ;
        RECT 134.00 19.00 141.00 21.00 ;
        RECT 14.00 19.00 46.00 21.00 ;
        RECT 29.00 24.00 52.00 26.00 ;
        RECT 19.00 24.00 26.00 26.00 ;
        RECT 62.00 19.00 76.00 21.00 ;
        RECT 86.00 24.00 100.00 26.00 ;
        RECT 110.00 19.00 124.00 21.00 ;
        RECT 134.00 24.00 148.00 26.00 ;
        RECT 19.00 24.00 151.00 26.00 ;
        LAYER L_ALU3 ;
        RECT 119.00 -1.00 131.00 51.00 ;
        RECT -6.00 -1.00 6.00 51.00 ;
    END
END ram_sense_buf0


MACRO ram_sense_buf1
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      170.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nwrite
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 94.00 29.00 96.00 31.00 ;
        END
    END nwrite
    PIN nckx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 104.00 29.00 106.00 31.00 ;
        END
    END nckx
    PIN nsense
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 69.00 29.00 71.00 31.00 ;
        END
    END nsense
    PIN selramx
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 54.00 29.00 56.00 31.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 34.00 29.00 36.00 31.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 24.00 29.00 26.00 31.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END selramx
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 154.00 24.00 156.00 26.00 ;
            RECT 149.00 24.00 151.00 26.00 ;
            RECT 144.00 24.00 146.00 26.00 ;
            RECT 139.00 24.00 141.00 26.00 ;
            RECT 134.00 24.00 136.00 26.00 ;
            RECT 129.00 24.00 131.00 26.00 ;
            RECT 124.00 24.00 126.00 26.00 ;
            RECT 119.00 24.00 121.00 26.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
            RECT 109.00 24.00 111.00 26.00 ;
            RECT 104.00 24.00 106.00 26.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 94.00 24.00 96.00 26.00 ;
            RECT 89.00 24.00 91.00 26.00 ;
            RECT 84.00 24.00 86.00 26.00 ;
            RECT 79.00 24.00 81.00 26.00 ;
            RECT 74.00 24.00 76.00 26.00 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 64.00 24.00 66.00 26.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
        END
    END nck
    PIN w
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 84.00 34.00 86.00 36.00 ;
            RECT 84.00 29.00 86.00 31.00 ;
            RECT 84.00 24.00 86.00 26.00 ;
            RECT 84.00 19.00 86.00 21.00 ;
            RECT 84.00 14.00 86.00 16.00 ;
        END
    END w
    PIN selram
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END selram
    PIN ck
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 159.00 39.00 161.00 41.00 ;
            RECT 159.00 34.00 161.00 36.00 ;
            RECT 159.00 29.00 161.00 31.00 ;
            RECT 159.00 24.00 161.00 26.00 ;
            RECT 159.00 19.00 161.00 21.00 ;
            RECT 159.00 14.00 161.00 16.00 ;
            RECT 159.00 9.00 161.00 11.00 ;
        END
    END ck
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 167.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 167.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 168.50 41.00 ;
        LAYER L_ALU2 ;
        RECT -1.00 -6.00 131.00 6.00 ;
        RECT -1.00 44.00 131.00 56.00 ;
        RECT 69.00 29.00 76.00 31.00 ;
        RECT 104.00 29.00 111.00 31.00 ;
        RECT 69.00 29.00 111.00 31.00 ;
        RECT 89.00 29.00 96.00 31.00 ;
        LAYER L_ALU3 ;
        RECT 119.00 -1.00 131.00 51.00 ;
        RECT -6.00 -1.00 6.00 51.00 ;
    END
END ram_sense_buf1


MACRO ram_sense_data
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      170.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN dout
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 99.00 39.00 101.00 41.00 ;
            RECT 99.00 34.00 101.00 36.00 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 99.00 24.00 101.00 26.00 ;
            RECT 99.00 19.00 101.00 21.00 ;
            RECT 99.00 14.00 101.00 16.00 ;
            RECT 99.00 9.00 101.00 11.00 ;
        END
    END dout
    PIN din
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 164.00 34.00 166.00 36.00 ;
            RECT 164.00 29.00 166.00 31.00 ;
            RECT 164.00 24.00 166.00 26.00 ;
            RECT 164.00 19.00 166.00 21.00 ;
        END
    END din
    PIN prechx
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 39.00 116.00 41.00 ;
            RECT 114.00 34.00 116.00 36.00 ;
            RECT 114.00 29.00 116.00 31.00 ;
            RECT 114.00 24.00 116.00 26.00 ;
            RECT 114.00 19.00 116.00 21.00 ;
            RECT 114.00 14.00 116.00 16.00 ;
            RECT 114.00 9.00 116.00 11.00 ;
        END
    END prechx
    PIN writex
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 134.00 34.00 136.00 36.00 ;
            RECT 134.00 29.00 136.00 31.00 ;
            RECT 134.00 24.00 136.00 26.00 ;
            RECT 134.00 19.00 136.00 21.00 ;
            RECT 134.00 14.00 136.00 16.00 ;
        END
    END writex
    PIN sensex
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 74.00 19.00 76.00 21.00 ;
        END
    END sensex
    PIN nsensex
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 24.00 91.00 26.00 ;
        END
    END nsensex
    PIN nbit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 39.00 26.00 41.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 9.00 39.00 11.00 41.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT -1.00 39.00 1.00 41.00 ;
        END
    END nbit1
    PIN bit1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 9.00 29.00 11.00 31.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT -1.00 29.00 1.00 31.00 ;
        END
    END bit1
    PIN bit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 24.00 9.00 26.00 11.00 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
            RECT -1.00 9.00 1.00 11.00 ;
        END
    END bit0
    PIN nbit0
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 9.00 19.00 11.00 21.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT -1.00 19.00 1.00 21.00 ;
        END
    END nbit0
    PIN nad0x
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END nad0x
    PIN ad0x
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END ad0x
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 167.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 167.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 168.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 89.00 24.00 161.00 26.00 ;
        RECT 146.00 24.00 161.00 26.00 ;
        RECT 118.00 39.00 155.00 41.00 ;
        RECT 89.00 39.00 155.00 41.00 ;
        RECT 89.00 9.00 143.00 11.00 ;
        RECT 118.00 9.00 143.00 11.00 ;
        RECT 56.00 19.00 81.00 21.00 ;
        RECT 29.00 19.00 36.00 21.00 ;
        RECT 29.00 39.00 36.00 41.00 ;
        RECT 84.00 24.00 91.00 26.00 ;
        RECT 19.00 21.00 21.00 31.00 ;
        RECT -1.00 9.00 91.00 41.00 ;
        RECT 10.00 34.00 16.00 36.00 ;
        RECT 10.00 14.00 16.00 16.00 ;
        RECT 134.00 14.00 141.00 16.00 ;
        RECT 134.00 34.00 141.00 36.00 ;
        RECT 89.00 34.00 141.00 36.00 ;
        RECT 89.00 14.00 141.00 16.00 ;
        RECT 19.00 34.00 125.00 36.00 ;
        RECT 19.00 14.00 125.00 16.00 ;
        RECT 109.00 24.00 116.00 26.00 ;
        LAYER L_ALU3 ;
        RECT -6.00 -1.00 6.00 51.00 ;
        RECT 119.00 -1.00 131.00 51.00 ;
    END
END ram_sense_data


MACRO ram_sense_decad12
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      170.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN ndec11
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 99.00 29.00 101.00 31.00 ;
            RECT 94.00 29.00 96.00 31.00 ;
        END
    END ndec11
    PIN ndec10
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 69.00 24.00 71.00 26.00 ;
            RECT 64.00 24.00 66.00 26.00 ;
        END
    END ndec10
    PIN ndec01
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END ndec01
    PIN ndec00
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END ndec00
    PIN ad2
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 139.00 39.00 141.00 41.00 ;
            RECT 139.00 34.00 141.00 36.00 ;
            RECT 139.00 29.00 141.00 31.00 ;
            RECT 139.00 24.00 141.00 26.00 ;
            RECT 139.00 19.00 141.00 21.00 ;
            RECT 139.00 14.00 141.00 16.00 ;
            RECT 139.00 9.00 141.00 11.00 ;
        END
    END ad2
    PIN ad1
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU1 ;
            RECT 164.00 39.00 166.00 41.00 ;
            RECT 164.00 34.00 166.00 36.00 ;
            RECT 164.00 29.00 166.00 31.00 ;
            RECT 164.00 24.00 166.00 26.00 ;
            RECT 164.00 19.00 166.00 21.00 ;
            RECT 164.00 14.00 166.00 16.00 ;
            RECT 164.00 9.00 166.00 11.00 ;
        END
    END ad1
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 167.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 167.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 168.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 76.00 9.00 146.00 11.00 ;
        RECT 16.00 14.00 141.00 16.00 ;
        RECT 22.00 39.00 166.00 41.00 ;
        RECT 52.00 34.00 161.00 36.00 ;
        RECT 22.00 39.00 166.00 41.00 ;
        RECT 52.00 34.00 161.00 36.00 ;
        RECT 16.00 14.00 141.00 16.00 ;
        RECT 76.00 9.00 146.00 11.00 ;
        LAYER L_ALU3 ;
        RECT -6.00 -1.00 6.00 51.00 ;
        RECT 119.00 -1.00 131.00 51.00 ;
    END
END ram_sense_decad12


MACRO ram_sense_decad2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      170.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN ad3x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 139.00 19.00 141.00 21.00 ;
        END
    END ad3x
    PIN nad3x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 154.00 19.00 156.00 21.00 ;
        END
    END nad3x
    PIN nad4x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 19.00 116.00 21.00 ;
        END
    END nad4x
    PIN ad4x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 19.00 111.00 21.00 ;
        END
    END ad4x
    PIN ad4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 134.00 19.00 136.00 21.00 ;
        END
    END ad4
    PIN ad3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 164.00 19.00 166.00 21.00 ;
        END
    END ad3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 167.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 167.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 168.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 104.00 19.00 166.00 21.00 ;
        RECT 139.00 19.00 146.00 21.00 ;
        RECT 159.00 19.00 166.00 21.00 ;
        RECT 149.00 19.00 156.00 21.00 ;
        RECT 129.00 19.00 136.00 21.00 ;
        RECT 104.00 19.00 111.00 21.00 ;
        RECT 114.00 19.00 123.00 21.00 ;
        LAYER L_ALU3 ;
        RECT -6.00 -1.00 6.00 51.00 ;
        RECT 119.00 -1.00 131.00 51.00 ;
    END
END ram_sense_decad2


MACRO ram_sense_decad3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      170.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nad5x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 19.00 91.00 21.00 ;
        END
    END nad5x
    PIN ad5x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 19.00 81.00 21.00 ;
        END
    END ad5x
    PIN ad3x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 139.00 19.00 141.00 21.00 ;
        END
    END ad3x
    PIN nad3x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 154.00 19.00 156.00 21.00 ;
        END
    END nad3x
    PIN nad4x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 19.00 116.00 21.00 ;
        END
    END nad4x
    PIN ad4x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 19.00 111.00 21.00 ;
        END
    END ad4x
    PIN ad5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 19.00 101.00 21.00 ;
        END
    END ad5
    PIN ad4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 134.00 19.00 136.00 21.00 ;
        END
    END ad4
    PIN ad3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 164.00 19.00 166.00 21.00 ;
        END
    END ad3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 167.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 167.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 168.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 74.00 19.00 166.00 21.00 ;
        RECT 104.00 19.00 111.00 21.00 ;
        RECT 94.00 19.00 101.00 21.00 ;
        RECT 84.00 19.00 91.00 21.00 ;
        RECT 74.00 19.00 81.00 21.00 ;
        RECT 129.00 19.00 136.00 21.00 ;
        RECT 139.00 19.00 146.00 21.00 ;
        RECT 149.00 19.00 156.00 21.00 ;
        RECT 159.00 19.00 166.00 21.00 ;
        RECT 114.00 19.00 123.00 21.00 ;
        LAYER L_ALU3 ;
        RECT -6.00 -1.00 6.00 51.00 ;
        RECT 119.00 -1.00 131.00 51.00 ;
    END
END ram_sense_decad3


MACRO ram_sense_decad4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      170.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN ad6x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END ad6x
    PIN nad6x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 54.00 19.00 56.00 21.00 ;
        END
    END nad6x
    PIN nad5x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 19.00 91.00 21.00 ;
        END
    END nad5x
    PIN ad5x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 19.00 81.00 21.00 ;
        END
    END ad5x
    PIN ad3x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 139.00 19.00 141.00 21.00 ;
        END
    END ad3x
    PIN nad3x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 154.00 19.00 156.00 21.00 ;
        END
    END nad3x
    PIN nad4x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 19.00 116.00 21.00 ;
        END
    END nad4x
    PIN ad4x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 19.00 111.00 21.00 ;
        END
    END ad4x
    PIN ad5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 19.00 101.00 21.00 ;
        END
    END ad5
    PIN ad6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 19.00 66.00 21.00 ;
        END
    END ad6
    PIN ad4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 134.00 19.00 136.00 21.00 ;
        END
    END ad4
    PIN ad3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 164.00 19.00 166.00 21.00 ;
        END
    END ad3
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 167.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 167.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 168.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 159.00 19.00 166.00 21.00 ;
        RECT 139.00 19.00 146.00 21.00 ;
        RECT 149.00 19.00 156.00 21.00 ;
        RECT 129.00 19.00 136.00 21.00 ;
        RECT 104.00 19.00 111.00 21.00 ;
        RECT 94.00 19.00 101.00 21.00 ;
        RECT 84.00 19.00 91.00 21.00 ;
        RECT 74.00 19.00 81.00 21.00 ;
        RECT 64.00 19.00 71.00 21.00 ;
        RECT 54.00 19.00 61.00 21.00 ;
        RECT 44.00 19.00 51.00 21.00 ;
        RECT 114.00 19.00 123.00 21.00 ;
        RECT 44.00 19.00 166.00 21.00 ;
        LAYER L_ALU3 ;
        RECT -6.00 -1.00 6.00 51.00 ;
        RECT 119.00 -1.00 131.00 51.00 ;
    END
END ram_sense_decad4


MACRO ram_sense_decad5
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      170.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN ad6x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END ad6x
    PIN nad6x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 54.00 19.00 56.00 21.00 ;
        END
    END nad6x
    PIN nad5x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 89.00 19.00 91.00 21.00 ;
        END
    END nad5x
    PIN ad5x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 79.00 19.00 81.00 21.00 ;
        END
    END ad5x
    PIN ad3x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 139.00 19.00 141.00 21.00 ;
        END
    END ad3x
    PIN nad3x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 154.00 19.00 156.00 21.00 ;
        END
    END nad3x
    PIN nad4x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 114.00 19.00 116.00 21.00 ;
        END
    END nad4x
    PIN ad7x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END ad7x
    PIN nad7x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END nad7x
    PIN ad4x
        DIRECTION OUTPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 109.00 19.00 111.00 21.00 ;
        END
    END ad4x
    PIN ad5
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 99.00 19.00 101.00 21.00 ;
        END
    END ad5
    PIN ad6
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 64.00 19.00 66.00 21.00 ;
        END
    END ad6
    PIN ad4
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 134.00 19.00 136.00 21.00 ;
        END
    END ad4
    PIN ad3
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 164.00 19.00 166.00 21.00 ;
        END
    END ad3
    PIN ad7
        DIRECTION INPUT ;
        PORT
            LAYER L_ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END ad7
    PIN vdd
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 167.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
            LAYER L_ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 167.00 3.00 ;
        END
    END vss
    OBS
        LAYER L_ALU1 ;
        RECT 1.50 9.00 168.50 41.00 ;
        LAYER L_ALU2 ;
        RECT 114.00 19.00 123.00 21.00 ;
        RECT 14.00 19.00 166.00 21.00 ;
        RECT 14.00 19.00 21.00 21.00 ;
        RECT 24.00 19.00 31.00 21.00 ;
        RECT 44.00 19.00 51.00 21.00 ;
        RECT 54.00 19.00 61.00 21.00 ;
        RECT 64.00 19.00 71.00 21.00 ;
        RECT 34.00 19.00 41.00 21.00 ;
        RECT 74.00 19.00 81.00 21.00 ;
        RECT 84.00 19.00 91.00 21.00 ;
        RECT 94.00 19.00 101.00 21.00 ;
        RECT 104.00 19.00 111.00 21.00 ;
        RECT 129.00 19.00 136.00 21.00 ;
        RECT 159.00 19.00 166.00 21.00 ;
        RECT 149.00 19.00 156.00 21.00 ;
        RECT 139.00 19.00 146.00 21.00 ;
        LAYER L_ALU3 ;
        RECT 119.00 -1.00 131.00 51.00 ;
        RECT -6.00 -1.00 6.00 51.00 ;
    END
END ram_sense_decad5


END LIBRARY
